  parameter integer NInstructions = 9;

  task startTest();                                                             // Free: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   2] = 'b0000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // free
      code[   3] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   4] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   5] = 'b0000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // free
      code[   6] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   7] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   8] = 'b0000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000001000000100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // free
    end
  endtask

  task endTest();                                                               // Free: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 0;
      success = success && outMem[1] == 0;
      success = success && outMem[2] == 0;
    end
  endtask
