  task startTest();                                                             // Array_scans: load code
    begin
      NInstructionEnd = 28;

      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;                                                                          // array
      code[   1] = 'h0000002300000000000000000000150000000000000a20000000000000000000;                                                                          // mov
      code[   2] = 'h0000002300000000000000000001150000000000001420000000000000000000;                                                                          // mov
      code[   3] = 'h0000002300000000000000000002150000000000001e20000000000000000000;                                                                          // mov
      code[   4] = 'h00000005000000000000000000012100000000000000210000000000001e2000;                                                                          // arrayIndex
      code[   5] = 'h0000002700000000000000000000010000000000000121000000000000000000;                                                                          // out
      code[   6] = 'h0000000500000000000000000002210000000000000021000000000000142000;                                                                          // arrayIndex
      code[   7] = 'h0000002700000000000000000000010000000000000221000000000000000000;                                                                          // out
      code[   8] = 'h00000005000000000000000000032100000000000000210000000000000a2000;                                                                          // arrayIndex
      code[   9] = 'h0000002700000000000000000000010000000000000321000000000000000000;                                                                          // out
      code[  10] = 'h00000005000000000000000000042100000000000000210000000000000f2000;                                                                          // arrayIndex
      code[  11] = 'h0000002700000000000000000000010000000000000421000000000000000000;                                                                          // out
      code[  12] = 'h0000000300000000000000000005210000000000000021000000000000232000;                                                                          // arrayCountLess
      code[  13] = 'h0000002700000000000000000000010000000000000521000000000000000000;                                                                          // out
      code[  14] = 'h0000000300000000000000000006210000000000000021000000000000192000;                                                                          // arrayCountLess
      code[  15] = 'h0000002700000000000000000000010000000000000621000000000000000000;                                                                          // out
      code[  16] = 'h00000003000000000000000000072100000000000000210000000000000f2000;                                                                          // arrayCountLess
      code[  17] = 'h0000002700000000000000000000010000000000000721000000000000000000;                                                                          // out
      code[  18] = 'h0000000300000000000000000008210000000000000021000000000000052000;                                                                          // arrayCountLess
      code[  19] = 'h0000002700000000000000000000010000000000000821000000000000000000;                                                                          // out
      code[  20] = 'h0000000200000000000000000009210000000000000021000000000000232000;                                                                          // arrayCountGreater
      code[  21] = 'h0000002700000000000000000000010000000000000921000000000000000000;                                                                          // out
      code[  22] = 'h000000020000000000000000000a210000000000000021000000000000192000;                                                                          // arrayCountGreater
      code[  23] = 'h0000002700000000000000000000010000000000000a21000000000000000000;                                                                          // out
      code[  24] = 'h000000020000000000000000000b2100000000000000210000000000000f2000;                                                                          // arrayCountGreater
      code[  25] = 'h0000002700000000000000000000010000000000000b21000000000000000000;                                                                          // out
      code[  26] = 'h000000020000000000000000000c210000000000000021000000000000052000;                                                                          // arrayCountGreater
      code[  27] = 'h0000002700000000000000000000010000000000000c21000000000000000000;                                                                          // out
    end
  endtask

  task endTest();                                                               // Array_scans: Evaluate results in out channel
    begin
      success = 1;

    end
  endtask
