  task startTest();                                                             // MoveLong_test: load code
    begin
      NInstructionEnd = 12;

      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;                                                                          // array
      code[   1] = 'h0000000100000000000000000001210000000000000420000000000000000000;                                                                          // array
      code[   2] = 'h0000002300000000000000000000150000000000000b20000000000000000000;                                                                          // mov
      code[   3] = 'h0000002300000000000000000001150000000000001620000000000000000000;                                                                          // mov
      code[   4] = 'h0000002300000000000000000002150000000000002120000000000000000000;                                                                          // mov
      code[   5] = 'h0000002300000000000000000003150000000000002c20000000000000000000;                                                                          // mov
      code[   6] = 'h0000002300000000000000000004150000000000003720000000000000000000;                                                                          // mov
      code[   7] = 'h0000002300000000000000010000150000000000004220000000000000000000;                                                                          // mov
      code[   8] = 'h0000002300000000000000010001150000000000004d20000000000000000000;                                                                          // mov
      code[   9] = 'h0000002300000000000000010002150000000000005820000000000000000000;                                                                          // mov
      code[  10] = 'h0000002300000000000000010003150000000000006320000000000000000000;                                                                          // mov
      code[  11] = 'h0000002400000000000000000001150000000001000115000000000000022000;                                                                          // moveLong
    end
  endtask

  task endTest();                                                               // MoveLong_test: Evaluate results in out channel
    begin
      success = 1;

    end
  endtask
