  parameter integer NInstructions = 3;

  task startTest();                                                             // Push_test: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000110000000000010000000000;                                          // push
      code[   2] = 'b0000000000000000000000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000110000000000010000000000;                                          // push
    end
  endtask

  task endTest();                                                               // Push_test: Evaluate results in out channel
    begin
      success = 1;
    end
  endtask
