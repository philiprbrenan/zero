  parameter integer NInstructions = 9;

  task startTest();                                                             // In_test: load code
    begin

      code[   0] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[   1] = 'b0000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // inSize
      code[   2] = 'b0000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011000000000000011000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jFalse
      code[   3] = 'b0000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // in
      code[   4] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   5] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   6] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[   7] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111100111110000000010000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[   8] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
    end
  endtask

  task endTest();                                                               // In_test: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 3;
      success = success && outMem[1] == 33;
      success = success && outMem[2] == 2;
      success = success && outMem[3] == 22;
      success = success && outMem[4] == 1;
      success = success && outMem[5] == 11;
    end
  endtask
