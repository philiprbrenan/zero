  task Add_test();
    begin                                                                       // Add_test
      NInstructionEnd = 2;

      code[   0] = 'h0000000000000000000000000000210000000000000320000000000000022000;                                                                          // add
      code[   1] = 'h0000002700000000000000000000010000000000000021000000000000000000;                                                                          // out
    end
  endtask
