//-----------------------------------------------------------------------------
// Fpga implementation and testing of NWay Trees
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga(input[1:0] in, output[1:0] out);                                    // Run test programs
  wire[1:0] in, out;                                                            // Input and output lines
  parameter integer NTestPrograms  =   18;                                      // Number of test programs to run
  parameter integer NTestsExpected =  118;                                      // Number of test passes expected
  parameter integer showInstructionDetails = 0;                                 // Show details of each instruction as it is executed

  parameter integer NSteps         = 2500;                                      // Maximum number of instruction executions
  parameter integer NInstructions  = 2000;                                      // Number of instruction slots in code memory
  parameter integer NArea          =   10;                                      // Size of each area on the heap
  parameter integer NArrays        = 1000;                                      // Amount of heap memory
  parameter integer NHeap          = NArea*NArrays;                             // Amount of heap memory
  parameter integer NLocal         = 1000;                                      // Size of local memory
  parameter integer NIn            = 1000;                                      // Size of input area
  parameter integer NOut           = 1000;                                      // Size of output area
  parameter integer NFreedArrays   = 1000;                                      // Size of output area
  parameter integer NMemoryPrintX  =   20;                                      // Width of memory to print
  parameter integer NMemoryPrintLines = 1;                                      // Number of lines of memory to print

  reg signed [255:0] code[NInstructions];                                       // Code memory
  reg signed [ 64:0] arraySizes[NArrays];                                       // Size of each array
  reg signed [ 64:0] heapMem [NHeap];                                           // Heap memory
  reg signed [ 64:0] localMem[NLocal];                                          // Local memory
  reg signed [ 64:0] inMem[NIn];                                                // Input channel
  reg signed [ 64:0] outMem[NOut];                                              // Out channel
  reg signed [ 64:0] freedArrays[NFreedArrays];                                 // Freed arrays list implemented as a stack
  reg signed [ 64:0] arrayShift[NArea];                                         // Array shift area

  integer signed nSteps;                                                        // Number of instructions executed
  integer signed NInstructionEnd;                                               // Limit of instructions for the current program
  integer signed  inMemPos;                                                     // Current position in input channel
  integer signed  inMemEnd;                                                     // End of input channel, this is the next element that would have been added.
  integer signed outMemPos;                                                     // Position in output channel
  integer signed result;                                                        // Result of an instruction execution
  integer signed allocs;                                                        // Maximum number of array allocations in use at any one time
  integer signed freedArraysTop;                                                // Position in freed arrays stack
  integer signed test;                                                          // Tests passed
  integer signed testsPassed;                                                   // Tests passed
  integer signed testsFailed;                                                   // Tests failed
  integer signed i, j, k, l, p, q;                                              // Useful integers

//Tests

  task ok(integer signed test, string name);                                    // Check a single test result
    begin
      if (test == 1) begin
        testsPassed++;
      end
      else begin
        $display("Assertion %s FAILED", name);
        printMemory();
        testsFailed++;
      end
    end
  endtask

  task loadCode();                                                              // Load code to be tested for test
    begin
      case(test)
        1: Mov_test();
        2: Add_test();
        3: Subtract_test();
        4: Not_test();
        5: Array_test();
        6: Array_scans();
        7: Free_test();
        8: ShiftLeft_test();
        9: ShiftRight_test();
       10: Jeq_test();
       11: Shift_up_test();
       12: Shift_up_test_2();
       13: Push_test();
       14: Pop_test();
       15: Bubble_sort();
       16: MoveLong_test();
       17: NWayTree_1();
       18: begin; inMemPos = 0; inMem[0] = 33; inMem[1] = 22; inMem[2] = 11; inMemEnd = 3; In_test(); end
      endcase

      case(test)                                                                // Initialize memory except in specific cases
        99:;
        default: initializeMemory();
      endcase
    end
  endtask

  task printMemory();                                                           // Print memory so we now what to chec
    begin
      $write("Local:");
      $write("      "); for(i = 0; i < NMemoryPrintX; ++i) $write(" %4d", i); $display("");
      for(j = 0; j < NLocal; j += NMemoryPrintX) begin
        if (j < NMemoryPrintLines) begin
          for(i = 0; i < NMemoryPrintX; ++i) begin
            $write(" %4d", localMem[j+i]);
          end
          $display("");
        end
      end
      $write("Heap: ");
      for(i = 0; i < NMemoryPrintX; ++i) begin
        $write(" %4d", heapMem[i]);
      end
      $display("");
    end
  endtask

  task printOut();                                                              // Print the output channel
    begin
      $display("Out %7d", outMemPos);
      $write("      "); for(i = 0; i < NMemoryPrintX; ++i) $write(" %4d", i); $display("");
      for(i = 0; i < outMemPos; ++i) begin
        $write(" %4d", outMem[i]);
      end
      $display("");
    end
  endtask

  task checkResults();                                                          // Check results of test
    begin
      case(test)
        1: ok(outMem[0] == 1, "Mov 1");                                         // 1
        2: ok(outMem[0] == 5, "Add 1");                                         // 1
        3: ok(outMem[0] == 2, "Subtract 1");                                    // 1
        4: begin                                                                // 3
          ok(outMem[0] == 3, "Not 1.1");
          ok(outMem[1] == 0, "Not 1.2");
          ok(outMem[2] == 1, "Not 1.3");
        end
        5: begin                                                                // 4 => 10
          ok(localMem[0] ==  0, "Array 1.1");
          ok( heapMem[0] == 11, "Array 1.2");
          ok( heapMem[1] == 22, "Array 1.3");
          ok( arraySizes[0] == 2, "Array 1.4");
        end
        6: begin                                                                // 12 => 22
          ok(outMem[0] == 3, "scan 1.1"); ok(outMem[1] == 2, "scan 1.2"); ok(outMem[ 2] == 1, "scan 1.3"); ok(outMem[ 3] == 0, "scan 1.4");
          ok(outMem[4] == 3, "scan 2.1"); ok(outMem[5] == 2, "scan 2.2"); ok(outMem[ 6] == 1, "scan 2.3"); ok(outMem[ 7] == 0, "scan 2.4");
          ok(outMem[8] == 0, "scan 3.1"); ok(outMem[9] == 1, "scan 3.2"); ok(outMem[10] == 2, "scan 3.3"); ok(outMem[11] == 3, "scan 3.4");
        end
        7: begin                                                                // 3    => 25
          ok(outMem[0] == 0, "Free 1"); ok(outMem[1] == 0, "Free 2"); ok(outMem[2] == 0, "Free 3");
        end
        8: begin
          ok(localMem[0] == 2, "ShiftLeft");                                    // 1
        end
        9: begin
          ok(localMem[0] == 2, "ShiftRight");                                   // 1
        end
       10: begin
          ok(outMem[0] == 111, "Jeq_test 1");                                   // 1
          ok(outMem[1] == 333, "Jeq_test 2");                                   // 1 => 29
        end
       11: begin
          ok(arraySizes[0] ==  4, "ShiftUp 1 length");                          // 5 => 34
          ok(heapMem[0]    == 99, "ShiftUp 1 new");
          ok(heapMem[1]    ==  0, "ShiftUp 1 0");
          ok(heapMem[2]    ==  1, "ShiftUp 1 1");
          ok(heapMem[3]    ==  2, "ShiftUp 1 2");
        end
       12: begin
          ok(arraySizes[0] ==  4, "ShiftUp 2 length");                          // 5 => 39
          ok(heapMem[0]    ==  0, "ShiftUp 2 new");
          ok(heapMem[1]    ==  1, "ShiftUp 2 0");
          ok(heapMem[2]    == 99, "ShiftUp 2 1");
          ok(heapMem[3]    ==  2, "ShiftUp 2 2");
        end
       13: begin
          ok(arraySizes[0] ==  2, "Push 1 length");                             // 3 => 42
          ok(heapMem[0]    ==  1, "Push 1 1");
          ok(heapMem[1]    ==  2, "Push 1 2");
        end
       14: begin
          ok(arraySizes[0] ==  0, "Pop 1 length");                              // 3 => 45
          ok(outMem[0]     ==  2, "Pop 1.1");
          ok(outMem[1]     ==  1, "Pop 1.2");
        end
       15: begin
          ok(arraySizes[0] ==  8, "Bubble Sort length");                        // 9 => 54
          ok(heapMem[0]    ==  11, "Bubble Sort 1");
          ok(heapMem[1]    ==  22, "Bubble Sort 2");
          ok(heapMem[2]    ==  33, "Bubble Sort 3");
          ok(heapMem[3]    ==  44, "Bubble Sort 4");
          ok(heapMem[4]    ==  55, "Bubble Sort 5");
          ok(heapMem[5]    ==  66, "Bubble Sort 6");
          ok(heapMem[6]    ==  77, "Bubble Sort 7");
          ok(heapMem[7]    ==  88, "Bubble Sort 8");
        end
       16: begin
          ok(arraySizes[0]  ==   5, "MoveLong Length aaa");                     // 11 => 65
          ok(arraySizes[1]  ==   4, "MoveLong Length bbb");
          ok(heapMem[0]     ==  11, "MoveLong 1");
          ok(heapMem[1]     ==  77, "MoveLong 2");
          ok(heapMem[2]     ==  88, "MoveLong 3");
          ok(heapMem[3]     ==  44, "MoveLong 4");
          ok(heapMem[4]     ==  55, "MoveLong 5");
          ok(heapMem[10]    ==  66, "MoveLong 6");
          ok(heapMem[11]    ==  77, "MoveLong 7");
          ok(heapMem[12]    ==  88, "MoveLong 8");
          ok(heapMem[13]    ==  99, "MoveLong 9");
        end
       17: begin
          ok(heapMem[ 00] == 6,  "NT100"); ok(heapMem[  1] ==  4,  "NT101"); ok(heapMem [02] == 3,  "NT102"); ok(heapMem [03] == 2, "NT103");
          ok(heapMem[ 20] == 2,  "NT120"); ok(heapMem[ 21] ==  1,  "NT121"); ok(heapMem [22] == 0,  "NT122"); ok(heapMem [23] == 0, "NT123");  ok(heapMem [24] ==  3, "NT124");  ok(heapMem [25] ==  4,  "NT125"); ok(heapMem [26] == 11, "NT126");
          ok(heapMem[ 30] == 2,  "NT130"); ok(heapMem[ 31] ==  4,  "NT131");
          ok(heapMem[ 50] == 2,  "NT150"); ok(heapMem[ 51] ==  2,  "NT151"); ok(heapMem [52] == 2,  "NT152"); ok(heapMem [53] == 0, "NT153");  ok(heapMem [54] ==  6, "NT154");  ok(heapMem [55] ==  7,  "NT155"); ok(heapMem [56] ==  0, "NT156");
          ok(heapMem[ 60] == 0,  "NT160"); ok(heapMem[ 61] ==  1,  "NT161");

          ok(heapMem[ 80] == 1,  "NT180"); ok(heapMem[ 81] ==  3,  "NT181"); ok(heapMem [82] == 2,  "NT182"); ok(heapMem [83] == 0, "NT183");  ok(heapMem [84] ==  9, "NT184");  ok(heapMem [85] == 10,  "NT185"); ok(heapMem [86] ==  0, "NT186");
          ok(heapMem[ 90] == 5,  "NT190");
          ok(heapMem[110] == 5, "NT1110"); ok(heapMem[111] == 12, "NT1111"); ok(heapMem[112] == 8, "NT1112");
          ok(heapMem[120] == 1, "NT1120"); ok(heapMem[121] ==  4, "NT1121"); ok(heapMem[122] == 2, "NT1122"); ok(heapMem[123] == 0, "NT1123"); ok(heapMem[124] == 13, "NT1124"); ok(heapMem[125] == 14, "NT1125"); ok(heapMem[126] ==  0, "NT1126");
          ok(heapMem[140] == 3, "NT1140");

          ok(outMem[0] == 0, "NT1 Out 0"); ok(outMem[1] == 1, "NT1 Out 1"); ok(outMem[2] == 2, "NT1 Out 2");
          ok(outMem[3] == 3, "NT1 Out 3"); ok(outMem[4] == 4, "NT1 Out 4"); ok(outMem[5] == 5, "NT1 Out 5");
        end
       18: begin
          ok(outMem[0] ==  3, "In1"); ok(outMem[1] == 33, "In2");
          ok(outMem[2] ==  2, "In3"); ok(outMem[3] == 22, "In4");
          ok(outMem[4] ==  1, "In5"); ok(outMem[5] == 11, "In6");
        end
      endcase
    end
  endtask

//Layout of each instruction

  integer ip = 0;                                                               // Instruction pointer
  integer r1, r2, r3, r4, r5, r6, r7, r8;                                       // Intermediate array results

  wire signed [255:0] instruction = code[ip];
  wire signed [31:0]  operator    = instruction[255:224];
  wire signed [63:0]  source2     = instruction[ 63:  0];
  wire signed [63:0]  source      = instruction[127: 64];
  wire signed [63:0]  target      = instruction[191:128];

  wire signed [31: 0] source2Area     = source2[63:32];                         // Source 2
  wire signed [15: 0] source2Address  = source2[31:16];
  wire signed [ 2: 0] source2Arena    = source2[13:12];
  wire signed [ 2: 0] source2DArea    = source2[11:10];
  wire signed [ 2: 0] source2DAddress = source2[ 9: 8];
  wire signed [ 7: 0] source2Delta    = source2[ 7: 0];
  wire signed [31: 0] source2Value    =                                         // Source 2 as value
    source2Arena      == 0 ? 0 :
    source2Arena      == 1 ?
     (                        source2DAddress == 0 ? source2Address :
      source2DArea    == 0 && source2DAddress == 1 ? heapMem [source2Delta + source2Area*NArea           + source2Address]           :
      source2DArea    == 0 && source2DAddress == 2 ? heapMem [source2Delta + source2Area*NArea           + localMem[source2Address]] :
      source2DArea    == 1 && source2DAddress == 1 ? heapMem [source2Delta + localMem[source2Area]*NArea + source2Address]           :
      source2DArea    == 1 && source2DAddress == 2 ? heapMem [source2Delta + localMem[source2Area]*NArea + localMem[source2Address]] : 0) :
    source2Arena      == 2 ?
     (source2DAddress == 0 ? source2Address :
      source2DAddress == 1 ? localMem[source2Delta + source2Address]           :
      source2DAddress == 2 ? localMem[source2Delta + localMem[source2Address]] : 0) : 0;

  wire signed [31: 0] source1Area     = source[63:32];                          // Source 1
  wire signed [15: 0] source1Address  = source[31:16];
  wire signed [ 2: 0] source1Arena    = source[13:12];
  wire signed [ 2: 0] source1DArea    = source[11:10];
  wire signed [ 2: 0] source1DAddress = source[ 9: 8];
  wire signed [ 7: 0] source1Delta    = source[ 7: 0];
  wire signed [31: 0] source1Value    =                                         // Source 1 as value
    source1Arena      == 0 ? 0 :
    source1Arena      == 1 ?
     (                        source1DAddress == 0 ? source1Address :
      source1DArea    == 0 && source1DAddress == 1 ? heapMem [source1Delta + source1Area*NArea           + source1Address]           :
      source1DArea    == 0 && source1DAddress == 2 ? heapMem [source1Delta + source1Area*NArea           + localMem[source1Address]] :
      source1DArea    == 1 && source1DAddress == 1 ? heapMem [source1Delta + localMem[source1Area]*NArea + source1Address]           :
      source1DArea    == 1 && source1DAddress == 2 ? heapMem [source1Delta + localMem[source1Area]*NArea + localMem[source1Address]] : 0) :
    source1Arena      == 2 ?
     (source1DAddress == 0 ? source1Address :
      source1DAddress == 1 ? localMem[source1Delta + source1Address]           :
      source1DAddress == 2 ? localMem[source1Delta + localMem[source1Address]] : 0) : 0;
  wire signed [31: 0] sourceLocation  =                                         // Source 1 as a location
    source1Arena      == 0 ? 0 :
    source1Arena      == 1 ?
     (                        source1DAddress == 0 ? source1Address :
      source1DArea    == 0 && source1DAddress == 1 ? source1Delta + source1Area*NArea           + source1Address           :
      source1DArea    == 0 && source1DAddress == 2 ? source1Delta + source1Area*NArea           + localMem[source1Address] :
      source1DArea    == 1 && source1DAddress == 1 ? source1Delta + localMem[source1Area]*NArea + source1Address           :
      source1DArea    == 1 && source1DAddress == 2 ? source1Delta + localMem[source1Area]*NArea + localMem[source1Address] : 0) :
    source1Arena      == 2 ?
     (source1DAddress == 0 ? source1Address :
      source1DAddress == 1 ? source1Delta + localMem[source1Address]           :
      source1DAddress == 2 ? source1Delta + localMem[localMem[source1Address]] : 0) : 0;

  wire signed [31: 0] targetArea      = target[63:32];                          // Target
  wire signed [15: 0] targetAddress   = target[31:16];
  wire signed [ 2: 0] targetArena     = target[13:12];
  wire signed [ 2: 0] targetDArea     = target[11:10];
  wire signed [ 2: 0] targetDAddress  = target[ 9: 8];
  wire signed [ 7: 0] targetDelta     = target[ 7: 0];
  wire signed [31: 0] targetLocation  =                                         // Target as a location
    targetArena      == 0 ? 0 :                                                 // Invalid
    targetArena      == 1 ?                                                     // Heap
     (targetDArea    == 0 && targetDAddress == 1 ? targetDelta + targetArea*NArea           + targetAddress           :
      targetDArea    == 0 && targetDAddress == 2 ? targetDelta + targetArea*NArea           + localMem[targetAddress] :
      targetDArea    == 1 && targetDAddress == 1 ? targetDelta + localMem[targetArea]*NArea + targetAddress           :
      targetDArea    == 1 && targetDAddress == 2 ? targetDelta + localMem[targetArea]*NArea + localMem[targetAddress] : 0) :
    targetArena      == 2 ?                                                     // Local
     (targetDAddress == 1 ?  targetDelta + targetAddress           :
      targetDAddress == 2 ?  targetDelta + localMem[targetAddress] : 0) : 0;

  wire signed [31: 0] targetIndex  =                                            // Target index within array
    targetArena      == 1 ?                                                     // Heap
     (targetDAddress == 1 ? targetDelta + targetAddress           :
      targetDAddress == 2 ? targetDelta + localMem[targetAddress] : 0)  : 0;

  wire signed [31: 0] targetLocationArea =                                      // Number of array containing target
      targetArena    == 1 && targetDArea == 0 ? targetArea :
      targetArena    == 1 && targetDArea == 1 ? localMem[targetArea]    : 0;

  wire signed [31: 0] targetValue    =                                          // Target as value
    targetArena      == 0 ? 0 :
    targetArena      == 1 ?
     (                       targetDAddress == 0 ? targetAddress :
      targetDArea    == 0 && targetDAddress == 1 ? heapMem [targetDelta + targetArea*NArea           + targetAddress]           :
      targetDArea    == 0 && targetDAddress == 2 ? heapMem [targetDelta + targetArea*NArea           + localMem[targetAddress]] :
      targetDArea    == 1 && targetDAddress == 1 ? heapMem [targetDelta + localMem[targetArea]*NArea + targetAddress]           :
      targetDArea    == 1 && targetDAddress == 2 ? heapMem [targetDelta + localMem[targetArea]*NArea + localMem[targetAddress]] : 0) :
    targetArena      == 2 ?
     (targetDAddress == 0 ? targetAddress :
      targetDAddress == 1 ? localMem[targetDelta + targetAddress]           :
      targetDAddress == 2 ? localMem[targetDelta + localMem[targetAddress]] : 0) : 0;

  task printInstruction();                                                      // Print an instruction
    begin;
      $display("targetAddress =%4x Area=%4x DAddress=%4x DArea=%4x Arena=%4x Delta=%4x Location=%4x value=%4x",
        targetAddress, targetArea, targetDAddress, targetDArea, targetArena, targetDelta, targetLocation, targetValue);

      $display("source1Address=%4x Area=%4x DAddress=%4x DArea=%4x Arena=%4x Delta=%4x Value   =%4x",
        source1Address, source1Area, source1DAddress, source1DArea, source1Arena, source1Delta, source1Value);

      $display("source2Address=%4x Area=%4x DAddress=%4x DArea=%4x Arena=%4x Delta=%4x Value   =%4x",
        source2Address, source2Area, source2DAddress, source2DArea, source2Arena, source2Delta, source2Value);
    end
  endtask

  task initializeMemory();                                                      // Initialize memory so we start in a known state
    begin;
      allocs         = 0;                                                       // Largest number of arrays in use at any one time so far
      freedArraysTop = 0;                                                       // Start freed arrays stack
      outMemPos      = 0;                                                       // Output channel position
      nSteps         = 1;                                                       // Number of instructions executed
      for(i = 0; i < NOut;    ++i)     outMem[i] = 'bx;                         // Reset the output channel
      for(i = 0; i < NHeap;   ++i)    heapMem[i] = 'bx;                         // Reset heap memory
      for(i = 0; i < NLocal;  ++i)   localMem[i] = 'bx;                         // Reset local memory
      for(i = 0; i < NArrays; ++i) arraySizes[i] =  0;                          // Set array sizes
    end
  endtask


// Execute each test progam

  initial begin                                                                 // Load, run confirm
    testsPassed = 0;                                                            // Passed tests
    testsFailed = 0;                                                            // Failed tests
    for(test = 1; test <= NTestPrograms; ++test) begin                          // Run the tests from bewest to oldest
      loadCode();
//if (test == 18) begin
      for(ip = 0; ip >= 0 && ip < NInstructionEnd; ++ip)                        // Each instruction
      begin
        #1;                                                                     // Let the ip update its assigns
        if (showInstructionDetails) printInstruction();                         // Print Instruction details
//Execute
        executeInstruction();

        if (nSteps++ > NSteps) begin                                            // Count instructions executed
          $display("Out of instructions after %d steps", NSteps);
          printMemory();
          $finish;
        end
      end
      $display("Test %4d, steps %8d", test, nSteps);
      checkResults();                                                           // Check results
//end
    end
    if (testsPassed > 0 && testsFailed > 0) begin
       $display("Passed %1d tests, FAILED %1d tests out of %d tests", testsPassed, testsFailed, NTestsExpected);
    end
    else if (testsFailed > 0) begin
       $display("FAILED %1d tests out of %1d tests", testsFailed, NTestsExpected);
    end
    else if (testsPassed > 0 && testsPassed != NTestsExpected) begin
       $display("Passed %1d tests out of %1d tests with no failures ", testsPassed, NTestsExpected);
    end
    else if (testsPassed == NTestsExpected) begin                               // Testing summary
       $display("All %1d tests passed successfully in %1d programs", NTestsExpected, NTestPrograms);
    end
    else begin
       $display("No tests run passed: %1d, failed: %1d, expected %1d, programs: %1d", testsPassed, testsFailed, NTestsExpected, NTestPrograms);
    end
    $finish;
  end

//Single instruction execution

  task executeInstruction();                                                    // Execute an instruction
    begin
      result = 'bx;
      case(operator)
         0: begin; add_instruction();                                       end // add_instruction
         1: begin; array_instruction();                                     end // array_instruction
         2: begin; arrayCountGreater_instruction();                         end // arrayCountGreater_instruction
         3: begin; arrayCountLess_instruction();                            end // arrayCountLess_instruction
         4: begin; arrayDump_instruction();                                 end // arrayDump_instruction
         5: begin; arrayIndex_instruction();                                end // arrayIndex_instruction
         6: begin; arraySize_instruction();                                 end // arraySize_instruction
         7: begin; assert_instruction();                                    end // assert_instruction
         8: begin; assertEq_instruction();                                  end // assertEq_instruction
         9: begin; assertFalse_instruction();                               end // assertFalse_instruction
        10: begin; assertGe_instruction();                                  end // assertGe_instruction
        11: begin; assertGt_instruction();                                  end // assertGt_instruction
        12: begin; assertLe_instruction();                                  end // assertLe_instruction
        13: begin; assertLt_instruction();                                  end // assertLt_instruction
        14: begin; assertNe_instruction();                                  end // assertNe_instruction
        15: begin; assertTrue_instruction();                                end // assertTrue_instruction
        16: begin; call_instruction();                                      end // call_instruction
        17: begin; confess_instruction();                                   end // confess_instruction
        18: begin; dump_instruction();                                      end // dump_instruction
        19: begin; free_instruction();                                      end // free_instruction
        20: begin; in_instruction();                                        end // in_instruction
        21: begin; inSize_instruction();                                    end // inSize_instruction
        22: begin; jEq_instruction();                                       end // jEq_instruction
        23: begin; jFalse_instruction();                                    end // jFalse_instruction
        24: begin; jGe_instruction();                                       end // jGe_instruction
        25: begin; jGt_instruction();                                       end // jGt_instruction
        26: begin; jLe_instruction();                                       end // jLe_instruction
        27: begin; jLt_instruction();                                       end // jLt_instruction
        28: begin; jNe_instruction();                                       end // jNe_instruction
        29: begin; jTrue_instruction();                                     end // jTrue_instruction
        30: begin; jmp_instruction();                                       end // jmp_instruction
        31: begin; label_instruction();                                     end // label_instruction
        32: begin; loadAddress_instruction();                               end // loadAddress_instruction
        33: begin; loadArea_instruction();                                  end // loadArea_instruction
        34: begin; mov_instruction();                                       end // mov_instruction
        35: begin; moveLong_instruction();                                  end // moveLong_instruction
        36: begin; nop_instruction();                                       end // nop_instruction
        37: begin; not_instruction();                                       end // not_instruction
        38: begin; out_instruction();                                       end // out_instruction
        39: begin; parallelContinue_instruction();                          end // parallelContinue_instruction
        40: begin; parallelStart_instruction();                             end // parallelStart_instruction
        41: begin; parallelStop_instruction();                              end // parallelStop_instruction
        42: begin; paramsGet_instruction();                                 end // paramsGet_instruction
        43: begin; paramsPut_instruction();                                 end // paramsPut_instruction
        44: begin; pop_instruction();                                       end // pop_instruction
        45: begin; push_instruction();                                      end // push_instruction
        46: begin; random_instruction();                                    end // random_instruction
        47: begin; randomSeed_instruction();                                end // randomSeed_instruction
        48: begin; resize_instruction();                                    end // resize_instruction
        49: begin; return_instruction();                                    end // return_instruction
        50: begin; returnGet_instruction();                                 end // returnGet_instruction
        51: begin; returnPut_instruction();                                 end // returnPut_instruction
        52: begin; shiftDown_instruction();                                 end // shiftDown_instruction
        53: begin; shiftLeft_instruction();                                 end // shiftLeft_instruction
        54: begin; shiftRight_instruction();                                end // shiftRight_instruction
        55: begin; shiftUp_instruction();                                   end // shiftUp_instruction
        56: begin; subtract_instruction();                                  end // subtract_instruction
        57: begin; tally_instruction();                                     end // tally_instruction
        58: begin; trace_instruction();                                     end // trace_instruction
        59: begin; traceLabels_instruction();                               end // traceLabels_instruction
        60: begin; watch_instruction();                                     end // watch_instruction
      endcase
    end
  endtask
  task arrayDump_instruction();
    begin                                                                       // arrayDump
     $display("arrayDump");
    end
  endtask
  task assert_instruction();
    begin                                                                       // assert
     $display("assert");
    end
  endtask
  task assertEq_instruction();
    begin                                                                       // assertEq
     $display("assertEq");
    end
  endtask
  task assertFalse_instruction();
    begin                                                                       // assertFalse
     $display("assertFalse");
    end
  endtask
  task assertGe_instruction();
    begin                                                                       // assertGe
     $display("assertGe");
    end
  endtask
  task assertGt_instruction();
    begin                                                                       // assertGt
     $display("assertGt");
    end
  endtask
  task assertLe_instruction();
    begin                                                                       // assertLe
     $display("assertLe");
    end
  endtask
  task assertLt_instruction();
    begin                                                                       // assertLt
     $display("assertLt");
    end
  endtask
  task assertNe_instruction();
    begin                                                                       // assertNe
    //$display("assertNe");
    end
  endtask
  task assertTrue_instruction();
    begin                                                                       // assertTrue
     $display("assertTrue");
    end
  endtask
  task call_instruction();
    begin                                                                       // call
     $display("call");
    end
  endtask
  task confess_instruction();
    begin                                                                       // confess
     $display("confess");
    end
  endtask
  task dump_instruction();
    begin                                                                       // dump
     $display("dump");
    end
  endtask
  task label_instruction();
    begin                                                                       // label
    end
  endtask
  task loadAddress_instruction();
    begin                                                                       // loadAddress
     $display("loadAddress");
    end
  endtask
  task loadArea_instruction();
    begin                                                                       // loadArea
     $display("loadArea");
    end
  endtask
  task nop_instruction();
    begin                                                                       // nop
     $display("nop");
    end
  endtask
  task parallelContinue_instruction();
    begin                                                                       // parallelContinue
    //$display("parallelContinue");
    end
  endtask
  task parallelStart_instruction();
    begin                                                                       // parallelStart
    //$display("parallelStart");
    end
  endtask
  task parallelStop_instruction();
    begin                                                                       // parallelStop
    // $display("parallelStop");
    end
  endtask
  task paramsGet_instruction();
    begin                                                                       // paramsGet
     $display("paramsGet");
    end
  endtask
  task paramsPut_instruction();
    begin                                                                       // paramsPut
     $display("paramsPut");
    end
  endtask
  task random_instruction();
    begin                                                                       // random
     $display("random");
    end
  endtask
  task randomSeed_instruction();
    begin                                                                       // randomSeed
     $display("randomSeed");
    end
  endtask
  task return_instruction();
    begin                                                                       // return
     $display("return");
    end
  endtask
  task returnGet_instruction();
    begin                                                                       // returnGet
     $display("returnGet");
    end
  endtask
  task returnPut_instruction();
    begin                                                                       // returnPut
     $display("returnPut");
    end
  endtask
  task shiftDown_instruction();
    begin                                                                       // shiftDown
     $display("shiftDown");
    end
  endtask
  task tally_instruction();
    begin                                                                       // tally
     $display("tally");
    end
  endtask
  task trace_instruction();
    begin                                                                       // trace
     $display("trace");
    end
  endtask
  task traceLabels_instruction();
    begin                                                                       // traceLabels
     $display("traceLabels");
    end
  endtask
  task watch_instruction();
    begin                                                                       // watch
     $display("watch");
    end
  endtask

//Programs to execute as tests
  task Mov_test();                                                              // Load program 'Mov_test' into code memory
    begin
      NInstructionEnd = 6;
      code[   0] = 'h0000002200000000000000000000210000000000000120000000000000000000;
      code[   1] = 'h0000002200000000000000000001210000000000000220000000000000000000;
      code[   2] = 'h0000002200000000000000000002210000000000000320000000000000000000;
      code[   3] = 'h0000002600000000000000000000010000000000000021000000000000000000;
      code[   4] = 'h0000002600000000000000000000010000000000000121000000000000000000;
      code[   5] = 'h0000002600000000000000000000010000000000000221000000000000000000;
    end
  endtask

  task Add_test();                                                              // Load program 'Add_test' into code memory    begin
    begin
      NInstructionEnd = 2;
      code[   0] = 'h0000000000000000000000000000210000000000000320000000000000022000;
      code[   1] = 'h0000002600000000000000000000010000000000000021000000000000000000;
    end
  endtask

  task Not_test();                                                              // Load program 'Not_test' into code memory
    begin
      NInstructionEnd = 6;
      code[   0] = 'h0000002200000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002500000000000000000001210000000000000021000000000000000000;
      code[   2] = 'h0000002500000000000000000002210000000000000121000000000000000000;
      code[   3] = 'h0000002600000000000000000000010000000000000021000000000000000000;
      code[   4] = 'h0000002600000000000000000000010000000000000121000000000000000000;
      code[   5] = 'h0000002600000000000000000000010000000000000221000000000000000000;
    end
  endtask

  task Subtract_test();                                                         // Load program 'Subtract_test' into code memory
    begin
      NInstructionEnd = 2;
      code[   0] = 'h0000003800000000000000000000210000000000000420000000000000022000;
      code[   1] = 'h0000002600000000000000000000010000000000000021000000000000000000;
    end
  endtask

  task Array_test();                                                            // Load program 'Array_test' into code memory
    begin
      NInstructionEnd = 3;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002200000000000000000000150000000000000b20000000000000000000;
      code[   2] = 'h0000002200000000000000000001150000000000001620000000000000000000;
    end
  endtask
                                                                                // Load program 'Array_scans' into code memory
  task Array_scans();
    begin
      NInstructionEnd = 28;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002200000000000000000000150000000000000a20000000000000000000;
      code[   2] = 'h0000002200000000000000000001150000000000001420000000000000000000;
      code[   3] = 'h0000002200000000000000000002150000000000001e20000000000000000000;
      code[   4] = 'h00000005000000000000000000012100000000000000210000000000001e2000;
      code[   5] = 'h0000002600000000000000000000010000000000000121000000000000000000;
      code[   6] = 'h0000000500000000000000000002210000000000000021000000000000142000;
      code[   7] = 'h0000002600000000000000000000010000000000000221000000000000000000;
      code[   8] = 'h00000005000000000000000000032100000000000000210000000000000a2000;
      code[   9] = 'h0000002600000000000000000000010000000000000321000000000000000000;
      code[  10] = 'h00000005000000000000000000042100000000000000210000000000000f2000;
      code[  11] = 'h0000002600000000000000000000010000000000000421000000000000000000;
      code[  12] = 'h0000000300000000000000000005210000000000000021000000000000232000;
      code[  13] = 'h0000002600000000000000000000010000000000000521000000000000000000;
      code[  14] = 'h0000000300000000000000000006210000000000000021000000000000192000;
      code[  15] = 'h0000002600000000000000000000010000000000000621000000000000000000;
      code[  16] = 'h00000003000000000000000000072100000000000000210000000000000f2000;
      code[  17] = 'h0000002600000000000000000000010000000000000721000000000000000000;
      code[  18] = 'h0000000300000000000000000008210000000000000021000000000000052000;
      code[  19] = 'h0000002600000000000000000000010000000000000821000000000000000000;
      code[  20] = 'h0000000200000000000000000009210000000000000021000000000000232000;
      code[  21] = 'h0000002600000000000000000000010000000000000921000000000000000000;
      code[  22] = 'h000000020000000000000000000a210000000000000021000000000000192000;
      code[  23] = 'h0000002600000000000000000000010000000000000a21000000000000000000;
      code[  24] = 'h000000020000000000000000000b2100000000000000210000000000000f2000;
      code[  25] = 'h0000002600000000000000000000010000000000000b21000000000000000000;
      code[  26] = 'h000000020000000000000000000c210000000000000021000000000000052000;
      code[  27] = 'h0000002600000000000000000000010000000000000c21000000000000000000;
    end
  endtask

  task Free_test();
    begin
      NInstructionEnd = 9;
      code[   0] = 'h0000000100000000000000000000217f000000000003207f000000000000007f;
      code[   1] = 'h0000002600000000000000000000017f000000000000217f000000000000007f;
      code[   2] = 'h0000001300000000000000000000217f000000000003207f000000000000007f;
      code[   3] = 'h0000000100000000000000000001217f000000000004207f000000000000007f;
      code[   4] = 'h0000002600000000000000000000017f000000000001217f000000000000007f;
      code[   5] = 'h0000001300000000000000000001217f000000000004207f000000000000007f;
      code[   6] = 'h0000000100000000000000000002217f000000000005207f000000000000007f;
      code[   7] = 'h0000002600000000000000000000017f000000000002217f000000000000007f;
      code[   8] = 'h0000001300000000000000000002217f000000000005207f000000000000007f;
    end
  endtask
                                                                                // Load program 'ShiftLeft_test' into code memory
  task ShiftLeft_test();
    begin
      NInstructionEnd = 3;
      code[   0] = 'h0000002200000000000000000000210000000000000120000000000000000000;
      code[   1] = 'h0000003500000000000000000000210000000000000021000000000000000000;
      code[   2] = 'h0000002600000000000000000000010000000000000021000000000000000000;
    end
  endtask
                                                                                // Load program 'ShiftRight_test' into code memory
  task ShiftRight_test();
    begin
      NInstructionEnd = 3;
      code[   0] = 'h0000002200000000000000000000210000000000000120000000000000000000;
      code[   1] = 'h0000003500000000000000000000210000000000000021000000000000000000;
      code[   2] = 'h0000002600000000000000000000010000000000000021000000000000000000;
    end
  endtask

  task Jeq_test();
    begin
      NInstructionEnd = 12;
      code[   0] = 'h0000001f00000000000000000000010000000000000120000000000000000000;
      code[   1] = 'h0000002200000000000000000000210000000000000120000000000000000000;
      code[   2] = 'h0000002200000000000000000001210000000000000220000000000000000000;
      code[   3] = 'h0000001600000000000000050002210000000000000021000000000000012100;
      code[   4] = 'h0000002600000000000000000000010000000000006f20000000000000000000;
      code[   5] = 'h0000001600000000000000030002210000000000000021000000000000002100;
      code[   6] = 'h000000260000000000000000000001000000000000de20000000000000000000;
      code[   7] = 'h0000001e00000000000000040004210000000000000000000000000000000000;
      code[   8] = 'h0000001f00000000000000000000010000000000000220000000000000000000;
      code[   9] = 'h0000002600000000000000000000010000000000014d20000000000000000000;
      code[  10] = 'h0000001f00000000000000000000010000000000000320000000000000000000;
      code[  11] = 'h0000001f00000000000000000000010000000000000420000000000000000000;
    end
  endtask
                                                                                // Load program 'Shift_up_test' into code memory
  task Shift_up_test();
    begin
      NInstructionEnd = 5;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002200000000000000000000150000000000000020000000000000000000;
      code[   2] = 'h0000002200000000000000000001150000000000000120000000000000000000;
      code[   3] = 'h0000002200000000000000000002150000000000000220000000000000000000;
      code[   4] = 'h0000003700000000000000000000150000000000006320000000000000000000;
    end
  endtask
                                                                                // Load program 'Shift_up_test_2' into code memory
  task Shift_up_test_2();
    begin
      NInstructionEnd = 5;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002200000000000000000000150000000000000020000000000000000000;
      code[   2] = 'h0000002200000000000000000001150000000000000120000000000000000000;
      code[   3] = 'h0000002200000000000000000002150000000000000220000000000000000000;
      code[   4] = 'h0000003700000000000000000002150000000000006320000000000000000000;
    end
  endtask

  task Push_test();
    begin
      NInstructionEnd = 3;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002d00000000000000000000210000000000000120000000000000032000;
      code[   2] = 'h0000002d00000000000000000000210000000000000220000000000000032000;
    end
  endtask

  task Pop_test();
    begin
      NInstructionEnd = 7;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002d00000000000000000000210000000000000120000000000000032000;
      code[   2] = 'h0000002d00000000000000000000210000000000000220000000000000032000;
      code[   3] = 'h0000002c00000000000000000001210000000000000021000000000000032000;
      code[   4] = 'h0000002c00000000000000000002210000000000000021000000000000032000;
      code[   5] = 'h0000002600000000000000000000010000000000000121000000000000000000;
      code[   6] = 'h0000002600000000000000000000010000000000000221000000000000000000;
    end
  endtask
                                                                                // Load program 'Bubble_sort' into code memory
  task Bubble_sort();
    begin
      NInstructionEnd = 44;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000002d00000000000000000000210000000000002120000000000000032000;
      code[   2] = 'h0000002d00000000000000000000210000000000000b20000000000000032000;
      code[   3] = 'h0000002d00000000000000000000210000000000001620000000000000032000;
      code[   4] = 'h0000002d00000000000000000000210000000000002c20000000000000032000;
      code[   5] = 'h0000002d00000000000000000000210000000000004d20000000000000032000;
      code[   6] = 'h0000002d00000000000000000000210000000000003720000000000000032000;
      code[   7] = 'h0000002d00000000000000000000210000000000004220000000000000032000;
      code[   8] = 'h0000002d00000000000000000000210000000000005820000000000000032000;
      code[   9] = 'h0000000600000000000000000001210000000000000021000000000000032000;
      code[  10] = 'h0000001f00000000000000000000010000000000000120000000000000000000;
      code[  11] = 'h0000002200000000000000000002210000000000000020000000000000000000;
      code[  12] = 'h0000001f00000000000000000000010000000000000220000000000000000000;
      code[  13] = 'h0000001800000000000000160004210000000000000221000000000000012100;
      code[  14] = 'h0000003800000000000000000003210000000000000121000000000000022100;
      code[  15] = 'h0000002200000000000000000004210000000000000020000000000000000000;
      code[  16] = 'h0000001f00000000000000000000010000000000000520000000000000000000;
      code[  17] = 'h0000002200000000000000000005210000000000000120000000000000000000;
      code[  18] = 'h0000001f00000000000000000000010000000000000620000000000000000000;
      code[  19] = 'h00000018000000000000000b0008210000000000000521000000000000032100;
      code[  20] = 'h0000002200000000000000000006210000000000000516000000000000000000;
      code[  21] = 'h0000002200000000000000000007210000000000000516ff0000000000000000;
      code[  22] = 'h0000001800000000000000040009210000000000000621000000000000072100;
      code[  23] = 'h000000220000000000000000000516ff00000000000621000000000000000000;
      code[  24] = 'h0000002200000000000000000005160000000000000721000000000000000000;
      code[  25] = 'h0000000000000000000000000004210000000000000421000000000000012000;
      code[  26] = 'h0000001f00000000000000000000010000000000000920000000000000000000;
      code[  27] = 'h0000001f00000000000000000000010000000000000720000000000000000000;
      code[  28] = 'h0000000000000000000000000005210000000000000521000000000000012000;
      code[  29] = 'h0000001e00000000fffffff50006210000000000000000000000000000000000;
      code[  30] = 'h0000001f00000000000000000000010000000000000820000000000000000000;
      code[  31] = 'h0000001700000000000000040004210000000000000421000000000000000000;
      code[  32] = 'h0000001f00000000000000000000010000000000000320000000000000000000;
      code[  33] = 'h0000000000000000000000000002210000000000000221000000000000012000;
      code[  34] = 'h0000001e00000000ffffffea0002210000000000000000000000000000000000;
      code[  35] = 'h0000001f00000000000000000000010000000000000420000000000000000000;
      code[  36] = 'h0000002600000000000000000000010000000000000015000000000000000000;
      code[  37] = 'h0000002600000000000000000000010000000000000115000000000000000000;
      code[  38] = 'h0000002600000000000000000000010000000000000215000000000000000000;
      code[  39] = 'h0000002600000000000000000000010000000000000315000000000000000000;
      code[  40] = 'h0000002600000000000000000000010000000000000415000000000000000000;
      code[  41] = 'h0000002600000000000000000000010000000000000515000000000000000000;
      code[  42] = 'h0000002600000000000000000000010000000000000615000000000000000000;
      code[  43] = 'h0000002600000000000000000000010000000000000715000000000000000000;
    end
  endtask

  task MoveLong_test();
    begin
      NInstructionEnd = 12;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;
      code[   1] = 'h0000000100000000000000000001210000000000000420000000000000000000;
      code[   2] = 'h0000002200000000000000000000150000000000000b20000000000000000000;
      code[   3] = 'h0000002200000000000000000001150000000000001620000000000000000000;
      code[   4] = 'h0000002200000000000000000002150000000000002120000000000000000000;
      code[   5] = 'h0000002200000000000000000003150000000000002c20000000000000000000;
      code[   6] = 'h0000002200000000000000000004150000000000003720000000000000000000;
      code[   7] = 'h0000002200000000000000010000150000000000004220000000000000000000;
      code[   8] = 'h0000002200000000000000010001150000000000004d20000000000000000000;
      code[   9] = 'h0000002200000000000000010002150000000000005820000000000000000000;
      code[  10] = 'h0000002200000000000000010003150000000000006320000000000000000000;
      code[  11] = 'h0000002300000000000000000001150000000001000115000000000000022000;
    end
  endtask

  task NWayTree_1();
    begin
      NInstructionEnd = 1655;
      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;                                                                          // array
      code[   1] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[   2] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[   3] = 'h0000002200000000000000000002150000000000000320000000000000000000;                                                                          // mov
      code[   4] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[   5] = 'h0000002200000000000000000001150000000000000020000000000000000000;                                                                          // mov
      code[   6] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[   7] = 'h0000002200000000000000000000150000000000000020000000000000000000;                                                                          // mov
      code[   8] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[   9] = 'h0000002200000000000000000003150000000000000020000000000000000000;                                                                          // mov
      code[  10] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[  11] = 'h0000001f00000000000000000000010000000000000120000000000000000000;                                                                          // label
      code[  12] = 'h0000003800000000000000000001210000000000000620000000000000012000;                                                                          // subtract
      code[  13] = 'h0000003800000000000000000002210000000000000121000000000000062000;                                                                          // subtract
      code[  14] = 'h0000001f00000000000000000000010000000000000220000000000000000000;                                                                          // label
      code[  15] = 'h0000001b00000000000005c60004210000000000000121000000000000002000;                                                                          // jLt
      code[  16] = 'h0000000100000000000000000003210000000000000420000000000000000000;                                                                          // array
      code[  17] = 'h0000001f00000000000000000000010000000000000520000000000000000000;                                                                          // label
      code[  18] = 'h0000002200000000000000000004210000000000000315000000000000000000;                                                                          // mov
      code[  19] = 'h0000001c00000000000000190009210000000000000421000000000000002000;                                                                          // jNe
      code[  20] = 'h0000000100000000000000000005210000000000000520000000000000000000;                                                                          // array
      code[  21] = 'h0000002200000000000000050000150000000000000120000000000000000000;                                                                          // mov
      code[  22] = 'h0000002200000000000000050002150000000000000020000000000000000000;                                                                          // mov
      code[  23] = 'h0000000100000000000000000006210000000000000620000000000000000000;                                                                          // array
      code[  24] = 'h0000002200000000000000050004150000000000000621000000000000000000;                                                                          // mov
      code[  25] = 'h0000000100000000000000000007210000000000000720000000000000000000;                                                                          // array
      code[  26] = 'h0000002200000000000000050005150000000000000721000000000000000000;                                                                          // mov
      code[  27] = 'h0000002200000000000000050006150000000000000020000000000000000000;                                                                          // mov
      code[  28] = 'h0000002200000000000000050003150000000000000021000000000000000000;                                                                          // mov
      code[  29] = 'h0000000000000000000000000001150000000000000115000000000000012000;                                                                          // add
      code[  30] = 'h0000002200000000000000050001150000000000000115000000000000000000;                                                                          // mov
      code[  31] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[  32] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  33] = 'h0000002200000000000000000008210000000005000415000000000000000000;                                                                          // mov
      code[  34] = 'h0000002200000000000000080000150000000000000121000000000000000000;                                                                          // mov
      code[  35] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  36] = 'h0000002200000000000000000003150000000000000521000000000000000000;                                                                          // mov
      code[  37] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  38] = 'h0000000000000000000000000000150000000000000015000000000000012000;                                                                          // add
      code[  39] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  40] = 'h0000002200000000000000000009210000000005000515000000000000000000;                                                                          // mov
      code[  41] = 'h0000002200000000000000090000150000000000000121000000000000000000;                                                                          // mov
      code[  42] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[  43] = 'h0000001e00000000000005a50008210000000000000000000000000000000000;                                                                          // jmp
      code[  44] = 'h0000001f00000000000000000000010000000000000920000000000000000000;                                                                          // label
      code[  45] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[  46] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  47] = 'h000000220000000000000000000a210000000000000215000000000000000000;                                                                          // mov
      code[  48] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  49] = 'h000000220000000000000000000b210000000004000015000000000000000000;                                                                          // mov
      code[  50] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[  51] = 'h00000018000000000000002f000a210000000000000b210000000000000a2100;                                                                          // jGe
      code[  52] = 'h000000220000000000000000000c210000000004000215000000000000000000;                                                                          // mov
      code[  53] = 'h0000001c000000000000002c000b210000000000000c21000000000000002000;                                                                          // jNe
      code[  54] = 'h000000250000000000000000000d210000000004000615000000000000000000;                                                                          // not
      code[  55] = 'h000000160000000000000029000c210000000000000d21000000000000002000;                                                                          // jEq
      code[  56] = 'h000000220000000000000000000e210000000004000415000000000000000000;                                                                          // mov
      code[  57] = 'h000000050000000000000000000f210000000000000e21000000000000012100;                                                                          // arrayIndex
      code[  58] = 'h000000160000000000000005000d210000000000000f21000000000000002000;                                                                          // jEq
      code[  59] = 'h000000380000000000000000000f210000000000000f21000000000000012000;                                                                          // subtract
      code[  60] = 'h0000002200000000000000000010210000000004000515000000000000000000;                                                                          // mov
      code[  61] = 'h000000220000000000000010000f160000000000000121000000000000000000;                                                                          // mov
      code[  62] = 'h0000001e00000000000005920008210000000000000000000000000000000000;                                                                          // jmp
      code[  63] = 'h0000001f00000000000000000000010000000000000d20000000000000000000;                                                                          // label
      code[  64] = 'h0000000200000000000000000011210000000000000e21000000000000012100;                                                                          // arrayCountGreater
      code[  65] = 'h0000001c000000000000000e000e210000000000001121000000000000002000;                                                                          // jNe
      code[  66] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[  67] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  68] = 'h0000002200000000000000000012210000000004000415000000000000000000;                                                                          // mov
      code[  69] = 'h000000220000000000000012000b160000000000000121000000000000000000;                                                                          // mov
      code[  70] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  71] = 'h0000000000000000000000000000150000000000000015000000000000012000;                                                                          // add
      code[  72] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  73] = 'h0000002200000000000000000013210000000004000515000000000000000000;                                                                          // mov
      code[  74] = 'h000000220000000000000013000b160000000000000121000000000000000000;                                                                          // mov
      code[  75] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  76] = 'h0000000000000000000000040000150000000000000b21000000000000012000;                                                                          // add
      code[  77] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[  78] = 'h0000001e00000000000005820008210000000000000000000000000000000000;                                                                          // jmp
      code[  79] = 'h0000001f00000000000000000000010000000000000e20000000000000000000;                                                                          // label
      code[  80] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[  81] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  82] = 'h0000000300000000000000000014210000000000000e21000000000000012100;                                                                          // arrayCountLess
      code[  83] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[  84] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  85] = 'h0000002200000000000000000015210000000004000515000000000000000000;                                                                          // mov
      code[  86] = 'h0000003700000000000000150014160000000000000121000000000000000000;                                                                          // shiftUp
      code[  87] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  88] = 'h0000002200000000000000000016210000000004000415000000000000000000;                                                                          // mov
      code[  89] = 'h0000003700000000000000160014160000000000000121000000000000000000;                                                                          // shiftUp
      code[  90] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[  91] = 'h0000000000000000000000040000150000000004000015000000000000012000;                                                                          // add
      code[  92] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[  93] = 'h0000000000000000000000000000150000000000000015000000000000012000;                                                                          // add
      code[  94] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[  95] = 'h0000001e00000000000005710008210000000000000000000000000000000000;                                                                          // jmp
      code[  96] = 'h0000001f00000000000000000000010000000000000c20000000000000000000;                                                                          // label
      code[  97] = 'h0000001f00000000000000000000010000000000000b20000000000000000000;                                                                          // label
      code[  98] = 'h0000001f00000000000000000000010000000000000a20000000000000000000;                                                                          // label
      code[  99] = 'h0000002200000000000000000017210000000000000315000000000000000000;                                                                          // mov
      code[ 100] = 'h0000001f00000000000000000000010000000000000f20000000000000000000;                                                                          // label
      code[ 101] = 'h0000002200000000000000000019210000000017000015000000000000000000;                                                                          // mov
      code[ 102] = 'h000000220000000000000000001a210000000017000315000000000000000000;                                                                          // mov
      code[ 103] = 'h000000220000000000000000001b21000000001a000215000000000000000000;                                                                          // mov
      code[ 104] = 'h0000001b000000000000013a00112100000000000019210000000000001b2100;                                                                          // jLt
      code[ 105] = 'h000000220000000000000000001c210000000000001b21000000000000000000;                                                                          // mov
      code[ 106] = 'h000000360000000000000000001c210000000000000120000000000000000000;                                                                          // shiftRight
      code[ 107] = 'h000000000000000000000000001d210000000000001c21000000000000012000;                                                                          // add
      code[ 108] = 'h000000220000000000000000001e210000000017000215000000000000000000;                                                                          // mov
      code[ 109] = 'h00000016000000000000008a0013210000000000001e21000000000000002000;                                                                          // jEq
      code[ 110] = 'h000000010000000000000000001f210000000000000520000000000000000000;                                                                          // array
      code[ 111] = 'h00000022000000000000001f0000150000000000001c21000000000000000000;                                                                          // mov
      code[ 112] = 'h00000022000000000000001f0002150000000000000020000000000000000000;                                                                          // mov
      code[ 113] = 'h0000000100000000000000000020210000000000000620000000000000000000;                                                                          // array
      code[ 114] = 'h00000022000000000000001f0004150000000000002021000000000000000000;                                                                          // mov
      code[ 115] = 'h0000000100000000000000000021210000000000000720000000000000000000;                                                                          // array
      code[ 116] = 'h00000022000000000000001f0005150000000000002121000000000000000000;                                                                          // mov
      code[ 117] = 'h00000022000000000000001f0006150000000000000020000000000000000000;                                                                          // mov
      code[ 118] = 'h00000022000000000000001f0003150000000000001a21000000000000000000;                                                                          // mov
      code[ 119] = 'h00000000000000000000001a000115000000001a000115000000000000012000;                                                                          // add
      code[ 120] = 'h00000022000000000000001f000115000000001a000115000000000000000000;                                                                          // mov
      code[ 121] = 'h0000002500000000000000000022210000000017000615000000000000000000;                                                                          // not
      code[ 122] = 'h0000001c00000000000000250014210000000000002221000000000000002000;                                                                          // jNe
      code[ 123] = 'h0000000100000000000000000023210000000000000820000000000000000000;                                                                          // array
      code[ 124] = 'h00000022000000000000001f0006150000000000002321000000000000000000;                                                                          // mov
      code[ 125] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 126] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 127] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 128] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 129] = 'h0000002200000000000000000024210000000017000515000000000000000000;                                                                          // mov
      code[ 130] = 'h000000220000000000000000002521000000001f000515000000000000000000;                                                                          // mov
      code[ 131] = 'h0000002300000000000000250000150000000024001d160000000000001c2100;                                                                          // moveLong
      code[ 132] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 133] = 'h0000002200000000000000000026210000000017000415000000000000000000;                                                                          // mov
      code[ 134] = 'h000000220000000000000000002721000000001f000415000000000000000000;                                                                          // mov
      code[ 135] = 'h0000002300000000000000270000150000000026001d160000000000001c2100;                                                                          // moveLong
      code[ 136] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 137] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 138] = 'h0000002200000000000000000028210000000017000615000000000000000000;                                                                          // mov
      code[ 139] = 'h000000220000000000000000002921000000001f000615000000000000000000;                                                                          // mov
      code[ 140] = 'h000000000000000000000000002a210000000000001c21000000000000012000;                                                                          // add
      code[ 141] = 'h0000002300000000000000290000150000000028001d160000000000002a2100;                                                                          // moveLong
      code[ 142] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 143] = 'h000000220000000000000000002b21000000001f000015000000000000000000;                                                                          // mov
      code[ 144] = 'h000000000000000000000000002c210000000000002b21000000000000012000;                                                                          // add
      code[ 145] = 'h000000220000000000000000002d21000000001f000615000000000000000000;                                                                          // mov
      code[ 146] = 'h0000001f00000000000000000000010000000000001620000000000000000000;                                                                          // label
      code[ 147] = 'h000000220000000000000000002e210000000000000020000000000000000000;                                                                          // mov
      code[ 148] = 'h0000001f00000000000000000000010000000000001720000000000000000000;                                                                          // label
      code[ 149] = 'h0000001800000000000000060019210000000000002e210000000000002c2100;                                                                          // jGe
      code[ 150] = 'h000000220000000000000000002f21000000002d002e16000000000000000000;                                                                          // mov
      code[ 151] = 'h00000022000000000000002f0002150000000000001f21000000000000000000;                                                                          // mov
      code[ 152] = 'h0000001f00000000000000000000010000000000001820000000000000000000;                                                                          // label
      code[ 153] = 'h000000000000000000000000002e210000000000002e21000000000000012000;                                                                          // add
      code[ 154] = 'h0000001e00000000fffffffa0017210000000000000000000000000000000000;                                                                          // jmp
      code[ 155] = 'h0000001f00000000000000000000010000000000001920000000000000000000;                                                                          // label
      code[ 156] = 'h0000002200000000000000000030210000000017000615000000000000000000;                                                                          // mov
      code[ 157] = 'h0000003000000000000000000030210000000000001d21000000000000082000;                                                                          // resize
      code[ 158] = 'h0000001e000000000000000c0015210000000000000000000000000000000000;                                                                          // jmp
      code[ 159] = 'h0000001f00000000000000000000010000000000001420000000000000000000;                                                                          // label
      code[ 160] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 161] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 162] = 'h0000002200000000000000000031210000000017000515000000000000000000;                                                                          // mov
      code[ 163] = 'h000000220000000000000000003221000000001f000515000000000000000000;                                                                          // mov
      code[ 164] = 'h0000002300000000000000320000150000000031001d160000000000001c2100;                                                                          // moveLong
      code[ 165] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 166] = 'h0000002200000000000000000033210000000017000415000000000000000000;                                                                          // mov
      code[ 167] = 'h000000220000000000000000003421000000001f000415000000000000000000;                                                                          // mov
      code[ 168] = 'h0000002300000000000000340000150000000033001d160000000000001c2100;                                                                          // moveLong
      code[ 169] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 170] = 'h0000001f00000000000000000000010000000000001520000000000000000000;                                                                          // label
      code[ 171] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 172] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 173] = 'h0000002200000000000000170000150000000000001c21000000000000000000;                                                                          // mov
      code[ 174] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 175] = 'h00000022000000000000001f0002150000000000001e21000000000000000000;                                                                          // mov
      code[ 176] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 177] = 'h000000220000000000000000003521000000001e000015000000000000000000;                                                                          // mov
      code[ 178] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 179] = 'h000000220000000000000000003621000000001e000615000000000000000000;                                                                          // mov
      code[ 180] = 'h0000002200000000000000000037210000000036003516000000000000000000;                                                                          // mov
      code[ 181] = 'h0000001c000000000000001c001a210000000000003721000000000000172100;                                                                          // jNe
      code[ 182] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 183] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 184] = 'h0000002200000000000000000038210000000017000515000000000000000000;                                                                          // mov
      code[ 185] = 'h0000002200000000000000000039210000000038001c16000000000000000000;                                                                          // mov
      code[ 186] = 'h000000220000000000000000003a21000000001e000515000000000000000000;                                                                          // mov
      code[ 187] = 'h00000022000000000000003a0035160000000000003921000000000000000000;                                                                          // mov
      code[ 188] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 189] = 'h000000220000000000000000003b210000000017000415000000000000000000;                                                                          // mov
      code[ 190] = 'h000000220000000000000000003c21000000003b001c16000000000000000000;                                                                          // mov
      code[ 191] = 'h000000220000000000000000003d21000000001e000415000000000000000000;                                                                          // mov
      code[ 192] = 'h00000022000000000000003d0035160000000000003c21000000000000000000;                                                                          // mov
      code[ 193] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 194] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 195] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 196] = 'h000000220000000000000000003e210000000017000515000000000000000000;                                                                          // mov
      code[ 197] = 'h000000300000000000000000003e210000000000001c21000000000000072000;                                                                          // resize
      code[ 198] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 199] = 'h000000220000000000000000003f210000000017000415000000000000000000;                                                                          // mov
      code[ 200] = 'h000000300000000000000000003f210000000000001c21000000000000062000;                                                                          // resize
      code[ 201] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 202] = 'h0000000000000000000000000040210000000000003521000000000000012000;                                                                          // add
      code[ 203] = 'h00000022000000000000001e0000150000000000004021000000000000000000;                                                                          // mov
      code[ 204] = 'h000000220000000000000000004121000000001e000615000000000000000000;                                                                          // mov
      code[ 205] = 'h0000002200000000000000410040160000000000001f21000000000000000000;                                                                          // mov
      code[ 206] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 207] = 'h0000001e00000000000000d00010210000000000000000000000000000000000;                                                                          // jmp
      code[ 208] = 'h0000001e0000000000000026001b210000000000000000000000000000000000;                                                                          // jmp
      code[ 209] = 'h0000001f00000000000000000000010000000000001a20000000000000000000;                                                                          // label
      code[ 210] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 211] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 212] = 'h0000000e00000000000000000000010000000000001e21000000000000002000;                                                                          // assertNe
      code[ 213] = 'h000000220000000000000000004221000000001e000615000000000000000000;                                                                          // mov
      code[ 214] = 'h0000000500000000000000000043210000000000004221000000000000172100;                                                                          // arrayIndex
      code[ 215] = 'h0000003800000000000000000043210000000000004321000000000000012000;                                                                          // subtract
      code[ 216] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 217] = 'h0000002200000000000000000044210000000017000415000000000000000000;                                                                          // mov
      code[ 218] = 'h0000002200000000000000000045210000000044001c16000000000000000000;                                                                          // mov
      code[ 219] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 220] = 'h0000002200000000000000000046210000000017000515000000000000000000;                                                                          // mov
      code[ 221] = 'h0000002200000000000000000047210000000046001c16000000000000000000;                                                                          // mov
      code[ 222] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 223] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 224] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 225] = 'h0000002200000000000000000048210000000017000515000000000000000000;                                                                          // mov
      code[ 226] = 'h0000003000000000000000000048210000000000001c21000000000000072000;                                                                          // resize
      code[ 227] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 228] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 229] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 230] = 'h000000220000000000000000004921000000001e000615000000000000000000;                                                                          // mov
      code[ 231] = 'h000000000000000000000000004a210000000000004321000000000000012000;                                                                          // add
      code[ 232] = 'h000000370000000000000049004a160000000000001f21000000000000000000;                                                                          // shiftUp
      code[ 233] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 234] = 'h000000220000000000000000004b21000000001e000415000000000000000000;                                                                          // mov
      code[ 235] = 'h00000037000000000000004b0043160000000000004521000000000000000000;                                                                          // shiftUp
      code[ 236] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 237] = 'h000000220000000000000000004c21000000001e000515000000000000000000;                                                                          // mov
      code[ 238] = 'h00000037000000000000004c0043160000000000004721000000000000000000;                                                                          // shiftUp
      code[ 239] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 240] = 'h00000000000000000000001e000015000000001e000015000000000000012000;                                                                          // add
      code[ 241] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 242] = 'h000000220000000000000000004d210000000017000415000000000000000000;                                                                          // mov
      code[ 243] = 'h000000300000000000000000004d210000000000001c21000000000000062000;                                                                          // resize
      code[ 244] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 245] = 'h0000001e00000000000000aa0010210000000000000000000000000000000000;                                                                          // jmp
      code[ 246] = 'h0000001f00000000000000000000010000000000001b20000000000000000000;                                                                          // label
      code[ 247] = 'h0000001f00000000000000000000010000000000001320000000000000000000;                                                                          // label
      code[ 248] = 'h000000010000000000000000004e210000000000000520000000000000000000;                                                                          // array
      code[ 249] = 'h00000022000000000000004e0000150000000000001c21000000000000000000;                                                                          // mov
      code[ 250] = 'h00000022000000000000004e0002150000000000000020000000000000000000;                                                                          // mov
      code[ 251] = 'h000000010000000000000000004f210000000000000620000000000000000000;                                                                          // array
      code[ 252] = 'h00000022000000000000004e0004150000000000004f21000000000000000000;                                                                          // mov
      code[ 253] = 'h0000000100000000000000000050210000000000000720000000000000000000;                                                                          // array
      code[ 254] = 'h00000022000000000000004e0005150000000000005021000000000000000000;                                                                          // mov
      code[ 255] = 'h00000022000000000000004e0006150000000000000020000000000000000000;                                                                          // mov
      code[ 256] = 'h00000022000000000000004e0003150000000000001a21000000000000000000;                                                                          // mov
      code[ 257] = 'h00000000000000000000001a000115000000001a000115000000000000012000;                                                                          // add
      code[ 258] = 'h00000022000000000000004e000115000000001a000115000000000000000000;                                                                          // mov
      code[ 259] = 'h0000000100000000000000000051210000000000000520000000000000000000;                                                                          // array
      code[ 260] = 'h0000002200000000000000510000150000000000001c21000000000000000000;                                                                          // mov
      code[ 261] = 'h0000002200000000000000510002150000000000000020000000000000000000;                                                                          // mov
      code[ 262] = 'h0000000100000000000000000052210000000000000620000000000000000000;                                                                          // array
      code[ 263] = 'h0000002200000000000000510004150000000000005221000000000000000000;                                                                          // mov
      code[ 264] = 'h0000000100000000000000000053210000000000000720000000000000000000;                                                                          // array
      code[ 265] = 'h0000002200000000000000510005150000000000005321000000000000000000;                                                                          // mov
      code[ 266] = 'h0000002200000000000000510006150000000000000020000000000000000000;                                                                          // mov
      code[ 267] = 'h0000002200000000000000510003150000000000001a21000000000000000000;                                                                          // mov
      code[ 268] = 'h00000000000000000000001a000115000000001a000115000000000000012000;                                                                          // add
      code[ 269] = 'h000000220000000000000051000115000000001a000115000000000000000000;                                                                          // mov
      code[ 270] = 'h0000002500000000000000000054210000000017000615000000000000000000;                                                                          // not
      code[ 271] = 'h0000001c000000000000004c001c210000000000005421000000000000002000;                                                                          // jNe
      code[ 272] = 'h0000000100000000000000000055210000000000000820000000000000000000;                                                                          // array
      code[ 273] = 'h00000022000000000000004e0006150000000000005521000000000000000000;                                                                          // mov
      code[ 274] = 'h0000000100000000000000000056210000000000000820000000000000000000;                                                                          // array
      code[ 275] = 'h0000002200000000000000510006150000000000005621000000000000000000;                                                                          // mov
      code[ 276] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 277] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 278] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 279] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 280] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 281] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 282] = 'h0000002200000000000000000057210000000017000415000000000000000000;                                                                          // mov
      code[ 283] = 'h0000002200000000000000000058210000000051000415000000000000000000;                                                                          // mov
      code[ 284] = 'h0000002300000000000000580000150000000057001d160000000000001c2100;                                                                          // moveLong
      code[ 285] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 286] = 'h0000002200000000000000000059210000000017000515000000000000000000;                                                                          // mov
      code[ 287] = 'h000000220000000000000000005a210000000051000515000000000000000000;                                                                          // mov
      code[ 288] = 'h00000023000000000000005a0000150000000059001d160000000000001c2100;                                                                          // moveLong
      code[ 289] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 290] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 291] = 'h000000220000000000000000005b210000000017000615000000000000000000;                                                                          // mov
      code[ 292] = 'h000000220000000000000000005c210000000051000615000000000000000000;                                                                          // mov
      code[ 293] = 'h000000000000000000000000005d210000000000001c21000000000000012000;                                                                          // add
      code[ 294] = 'h00000023000000000000005c000015000000005b001d160000000000005d2100;                                                                          // moveLong
      code[ 295] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 296] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 297] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 298] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 299] = 'h000000220000000000000000005e210000000017000615000000000000000000;                                                                          // mov
      code[ 300] = 'h000000220000000000000000005f21000000004e000615000000000000000000;                                                                          // mov
      code[ 301] = 'h0000000000000000000000000060210000000000001c21000000000000012000;                                                                          // add
      code[ 302] = 'h00000023000000000000005f000015000000005e000015000000000000602100;                                                                          // moveLong
      code[ 303] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 304] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 305] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 306] = 'h0000002200000000000000000061210000000017000415000000000000000000;                                                                          // mov
      code[ 307] = 'h000000220000000000000000006221000000004e000415000000000000000000;                                                                          // mov
      code[ 308] = 'h00000023000000000000006200001500000000610000150000000000001c2100;                                                                          // moveLong
      code[ 309] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 310] = 'h0000002200000000000000000063210000000017000515000000000000000000;                                                                          // mov
      code[ 311] = 'h000000220000000000000000006421000000004e000515000000000000000000;                                                                          // mov
      code[ 312] = 'h00000023000000000000006400001500000000630000150000000000001c2100;                                                                          // moveLong
      code[ 313] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 314] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 315] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 316] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 317] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 318] = 'h000000220000000000000000006521000000004e000015000000000000000000;                                                                          // mov
      code[ 319] = 'h0000000000000000000000000066210000000000006521000000000000012000;                                                                          // add
      code[ 320] = 'h000000220000000000000000006721000000004e000615000000000000000000;                                                                          // mov
      code[ 321] = 'h0000001f00000000000000000000010000000000001e20000000000000000000;                                                                          // label
      code[ 322] = 'h0000002200000000000000000068210000000000000020000000000000000000;                                                                          // mov
      code[ 323] = 'h0000001f00000000000000000000010000000000001f20000000000000000000;                                                                          // label
      code[ 324] = 'h0000001800000000000000060021210000000000006821000000000000662100;                                                                          // jGe
      code[ 325] = 'h0000002200000000000000000069210000000067006816000000000000000000;                                                                          // mov
      code[ 326] = 'h0000002200000000000000690002150000000000004e21000000000000000000;                                                                          // mov
      code[ 327] = 'h0000001f00000000000000000000010000000000002020000000000000000000;                                                                          // label
      code[ 328] = 'h0000000000000000000000000068210000000000006821000000000000012000;                                                                          // add
      code[ 329] = 'h0000001e00000000fffffffa001f210000000000000000000000000000000000;                                                                          // jmp
      code[ 330] = 'h0000001f00000000000000000000010000000000002120000000000000000000;                                                                          // label
      code[ 331] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 332] = 'h000000220000000000000000006a210000000051000015000000000000000000;                                                                          // mov
      code[ 333] = 'h000000000000000000000000006b210000000000006a21000000000000012000;                                                                          // add
      code[ 334] = 'h000000220000000000000000006c210000000051000615000000000000000000;                                                                          // mov
      code[ 335] = 'h0000001f00000000000000000000010000000000002220000000000000000000;                                                                          // label
      code[ 336] = 'h000000220000000000000000006d210000000000000020000000000000000000;                                                                          // mov
      code[ 337] = 'h0000001f00000000000000000000010000000000002320000000000000000000;                                                                          // label
      code[ 338] = 'h0000001800000000000000060025210000000000006d210000000000006b2100;                                                                          // jGe
      code[ 339] = 'h000000220000000000000000006e21000000006c006d16000000000000000000;                                                                          // mov
      code[ 340] = 'h00000022000000000000006e0002150000000000005121000000000000000000;                                                                          // mov
      code[ 341] = 'h0000001f00000000000000000000010000000000002420000000000000000000;                                                                          // label
      code[ 342] = 'h000000000000000000000000006d210000000000006d21000000000000012000;                                                                          // add
      code[ 343] = 'h0000001e00000000fffffffa0023210000000000000000000000000000000000;                                                                          // jmp
      code[ 344] = 'h0000001f00000000000000000000010000000000002520000000000000000000;                                                                          // label
      code[ 345] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 346] = 'h0000001e000000000000001d001d210000000000000000000000000000000000;                                                                          // jmp
      code[ 347] = 'h0000001f00000000000000000000010000000000001c20000000000000000000;                                                                          // label
      code[ 348] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 349] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 350] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 351] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 352] = 'h000000220000000000000000006f210000000017000415000000000000000000;                                                                          // mov
      code[ 353] = 'h000000220000000000000000007021000000004e000415000000000000000000;                                                                          // mov
      code[ 354] = 'h000000230000000000000070000015000000006f0000150000000000001c2100;                                                                          // moveLong
      code[ 355] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 356] = 'h0000002200000000000000000071210000000017000515000000000000000000;                                                                          // mov
      code[ 357] = 'h000000220000000000000000007221000000004e000515000000000000000000;                                                                          // mov
      code[ 358] = 'h00000023000000000000007200001500000000710000150000000000001c2100;                                                                          // moveLong
      code[ 359] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 360] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 361] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 362] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 363] = 'h0000002200000000000000000073210000000017000515000000000000000000;                                                                          // mov
      code[ 364] = 'h0000002200000000000000000074210000000051000515000000000000000000;                                                                          // mov
      code[ 365] = 'h0000002300000000000000740000150000000073001d160000000000001c2100;                                                                          // moveLong
      code[ 366] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 367] = 'h0000002200000000000000000075210000000017000415000000000000000000;                                                                          // mov
      code[ 368] = 'h0000002200000000000000000076210000000051000415000000000000000000;                                                                          // mov
      code[ 369] = 'h0000002300000000000000760000150000000075001d160000000000001c2100;                                                                          // moveLong
      code[ 370] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 371] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 372] = 'h0000000100000000000000000077210000000000000820000000000000000000;                                                                          // array
      code[ 373] = 'h0000002200000000000000170006150000000000007721000000000000000000;                                                                          // mov
      code[ 374] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 375] = 'h0000001f00000000000000000000010000000000001d20000000000000000000;                                                                          // label
      code[ 376] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 377] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 378] = 'h00000022000000000000004e0002150000000000001721000000000000000000;                                                                          // mov
      code[ 379] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 380] = 'h0000002200000000000000510002150000000000001721000000000000000000;                                                                          // mov
      code[ 381] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 382] = 'h0000002200000000000000000078210000000017000415000000000000000000;                                                                          // mov
      code[ 383] = 'h0000002200000000000000000079210000000078001c16000000000000000000;                                                                          // mov
      code[ 384] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 385] = 'h000000220000000000000000007a210000000017000515000000000000000000;                                                                          // mov
      code[ 386] = 'h000000220000000000000000007b21000000007a001c16000000000000000000;                                                                          // mov
      code[ 387] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 388] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 389] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 390] = 'h000000220000000000000000007c210000000017000615000000000000000000;                                                                          // mov
      code[ 391] = 'h00000022000000000000007c0001150000000000005121000000000000000000;                                                                          // mov
      code[ 392] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 393] = 'h000000220000000000000000007d210000000017000415000000000000000000;                                                                          // mov
      code[ 394] = 'h000000300000000000000000007d210000000000000120000000000000062000;                                                                          // resize
      code[ 395] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 396] = 'h000000220000000000000000007e210000000017000415000000000000000000;                                                                          // mov
      code[ 397] = 'h00000022000000000000007e0000150000000000007921000000000000000000;                                                                          // mov
      code[ 398] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 399] = 'h000000220000000000000000007f210000000017000515000000000000000000;                                                                          // mov
      code[ 400] = 'h00000022000000000000007f0000150000000000007b21000000000000000000;                                                                          // mov
      code[ 401] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 402] = 'h0000002200000000000000170000150000000000000120000000000000000000;                                                                          // mov
      code[ 403] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 404] = 'h0000002200000000000000000080210000000017000615000000000000000000;                                                                          // mov
      code[ 405] = 'h0000003000000000000000000080210000000000000220000000000000082000;                                                                          // resize
      code[ 406] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 407] = 'h0000002200000000000000000081210000000017000615000000000000000000;                                                                          // mov
      code[ 408] = 'h0000002200000000000000810000150000000000004e21000000000000000000;                                                                          // mov
      code[ 409] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 410] = 'h0000002200000000000000000082210000000017000515000000000000000000;                                                                          // mov
      code[ 411] = 'h0000003000000000000000000082210000000000000120000000000000072000;                                                                          // resize
      code[ 412] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 413] = 'h0000001e00000000000000020010210000000000000000000000000000000000;                                                                          // jmp
      code[ 414] = 'h0000001e00000000000000060012210000000000000000000000000000000000;                                                                          // jmp
      code[ 415] = 'h0000001f00000000000000000000010000000000001020000000000000000000;                                                                          // label
      code[ 416] = 'h0000002200000000000000000018210000000000000120000000000000000000;                                                                          // mov
      code[ 417] = 'h0000001e00000000000000030012210000000000000000000000000000000000;                                                                          // jmp
      code[ 418] = 'h0000001f00000000000000000000010000000000001120000000000000000000;                                                                          // label
      code[ 419] = 'h0000002200000000000000000018210000000000000020000000000000000000;                                                                          // mov
      code[ 420] = 'h0000001f00000000000000000000010000000000001220000000000000000000;                                                                          // label
      code[ 421] = 'h0000001f00000000000000000000010000000000002620000000000000000000;                                                                          // label
      code[ 422] = 'h0000001f00000000000000000000010000000000002a20000000000000000000;                                                                          // label
      code[ 423] = 'h0000002200000000000000000083210000000000000020000000000000000000;                                                                          // mov
      code[ 424] = 'h0000001f00000000000000000000010000000000002b20000000000000000000;                                                                          // label
      code[ 425] = 'h0000001800000000000002ba002d210000000000008321000000000000632000;                                                                          // jGe
      code[ 426] = 'h0000002200000000000000000084210000000017000015000000000000000000;                                                                          // mov
      code[ 427] = 'h0000003800000000000000000085210000000000008421000000000000012000;                                                                          // subtract
      code[ 428] = 'h0000002200000000000000000086210000000017000415000000000000000000;                                                                          // mov
      code[ 429] = 'h0000002200000000000000000087210000000086008516000000000000000000;                                                                          // mov
      code[ 430] = 'h0000001a0000000000000153002e210000000000000121000000000000872100;                                                                          // jLe
      code[ 431] = 'h0000002500000000000000000088210000000017000615000000000000000000;                                                                          // not
      code[ 432] = 'h000000160000000000000009002f210000000000008821000000000000002000;                                                                          // jEq
      code[ 433] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 434] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 435] = 'h0000002200000000000000030001150000000000000220000000000000000000;                                                                          // mov
      code[ 436] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 437] = 'h0000002200000000000000030000150000000000001721000000000000000000;                                                                          // mov
      code[ 438] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 439] = 'h0000003800000000000000030002150000000000008421000000000000012000;                                                                          // subtract
      code[ 440] = 'h0000001e00000000000002af0029210000000000000000000000000000000000;                                                                          // jmp
      code[ 441] = 'h0000001f00000000000000000000010000000000002f20000000000000000000;                                                                          // label
      code[ 442] = 'h0000002200000000000000000089210000000017000615000000000000000000;                                                                          // mov
      code[ 443] = 'h000000220000000000000000008a210000000089008416000000000000000000;                                                                          // mov
      code[ 444] = 'h0000001f00000000000000000000010000000000003020000000000000000000;                                                                          // label
      code[ 445] = 'h000000220000000000000000008c21000000008a000015000000000000000000;                                                                          // mov
      code[ 446] = 'h000000220000000000000000008d21000000008a000315000000000000000000;                                                                          // mov
      code[ 447] = 'h000000220000000000000000008e21000000008d000215000000000000000000;                                                                          // mov
      code[ 448] = 'h0000001b000000000000013a0032210000000000008c210000000000008e2100;                                                                          // jLt
      code[ 449] = 'h000000220000000000000000008f210000000000008e21000000000000000000;                                                                          // mov
      code[ 450] = 'h000000360000000000000000008f210000000000000120000000000000000000;                                                                          // shiftRight
      code[ 451] = 'h0000000000000000000000000090210000000000008f21000000000000012000;                                                                          // add
      code[ 452] = 'h000000220000000000000000009121000000008a000215000000000000000000;                                                                          // mov
      code[ 453] = 'h00000016000000000000008a0034210000000000009121000000000000002000;                                                                          // jEq
      code[ 454] = 'h0000000100000000000000000092210000000000000520000000000000000000;                                                                          // array
      code[ 455] = 'h0000002200000000000000920000150000000000008f21000000000000000000;                                                                          // mov
      code[ 456] = 'h0000002200000000000000920002150000000000000020000000000000000000;                                                                          // mov
      code[ 457] = 'h0000000100000000000000000093210000000000000620000000000000000000;                                                                          // array
      code[ 458] = 'h0000002200000000000000920004150000000000009321000000000000000000;                                                                          // mov
      code[ 459] = 'h0000000100000000000000000094210000000000000720000000000000000000;                                                                          // array
      code[ 460] = 'h0000002200000000000000920005150000000000009421000000000000000000;                                                                          // mov
      code[ 461] = 'h0000002200000000000000920006150000000000000020000000000000000000;                                                                          // mov
      code[ 462] = 'h0000002200000000000000920003150000000000008d21000000000000000000;                                                                          // mov
      code[ 463] = 'h00000000000000000000008d000115000000008d000115000000000000012000;                                                                          // add
      code[ 464] = 'h000000220000000000000092000115000000008d000115000000000000000000;                                                                          // mov
      code[ 465] = 'h000000250000000000000000009521000000008a000615000000000000000000;                                                                          // not
      code[ 466] = 'h0000001c00000000000000250035210000000000009521000000000000002000;                                                                          // jNe
      code[ 467] = 'h0000000100000000000000000096210000000000000820000000000000000000;                                                                          // array
      code[ 468] = 'h0000002200000000000000920006150000000000009621000000000000000000;                                                                          // mov
      code[ 469] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 470] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 471] = 'h000000220000000000000000009721000000008a000615000000000000000000;                                                                          // mov
      code[ 472] = 'h0000002200000000000000000098210000000092000615000000000000000000;                                                                          // mov
      code[ 473] = 'h0000000000000000000000000099210000000000008f21000000000000012000;                                                                          // add
      code[ 474] = 'h0000002300000000000000980000150000000097009016000000000000992100;                                                                          // moveLong
      code[ 475] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 476] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 477] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 478] = 'h000000220000000000000000009a21000000008a000415000000000000000000;                                                                          // mov
      code[ 479] = 'h000000220000000000000000009b210000000092000415000000000000000000;                                                                          // mov
      code[ 480] = 'h00000023000000000000009b000015000000009a0090160000000000008f2100;                                                                          // moveLong
      code[ 481] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 482] = 'h000000220000000000000000009c21000000008a000515000000000000000000;                                                                          // mov
      code[ 483] = 'h000000220000000000000000009d210000000092000515000000000000000000;                                                                          // mov
      code[ 484] = 'h00000023000000000000009d000015000000009c0090160000000000008f2100;                                                                          // moveLong
      code[ 485] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 486] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 487] = 'h000000220000000000000000009e210000000092000015000000000000000000;                                                                          // mov
      code[ 488] = 'h000000000000000000000000009f210000000000009e21000000000000012000;                                                                          // add
      code[ 489] = 'h00000022000000000000000000a0210000000092000615000000000000000000;                                                                          // mov
      code[ 490] = 'h0000001f00000000000000000000010000000000003720000000000000000000;                                                                          // label
      code[ 491] = 'h00000022000000000000000000a1210000000000000020000000000000000000;                                                                          // mov
      code[ 492] = 'h0000001f00000000000000000000010000000000003820000000000000000000;                                                                          // label
      code[ 493] = 'h000000180000000000000006003a21000000000000a1210000000000009f2100;                                                                          // jGe
      code[ 494] = 'h00000022000000000000000000a22100000000a000a116000000000000000000;                                                                          // mov
      code[ 495] = 'h0000002200000000000000a20002150000000000009221000000000000000000;                                                                          // mov
      code[ 496] = 'h0000001f00000000000000000000010000000000003920000000000000000000;                                                                          // label
      code[ 497] = 'h00000000000000000000000000a121000000000000a121000000000000012000;                                                                          // add
      code[ 498] = 'h0000001e00000000fffffffa0038210000000000000000000000000000000000;                                                                          // jmp
      code[ 499] = 'h0000001f00000000000000000000010000000000003a20000000000000000000;                                                                          // label
      code[ 500] = 'h00000022000000000000000000a321000000008a000615000000000000000000;                                                                          // mov
      code[ 501] = 'h00000030000000000000000000a3210000000000009021000000000000082000;                                                                          // resize
      code[ 502] = 'h0000001e000000000000000c0036210000000000000000000000000000000000;                                                                          // jmp
      code[ 503] = 'h0000001f00000000000000000000010000000000003520000000000000000000;                                                                          // label
      code[ 504] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 505] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 506] = 'h00000022000000000000000000a421000000008a000415000000000000000000;                                                                          // mov
      code[ 507] = 'h00000022000000000000000000a5210000000092000415000000000000000000;                                                                          // mov
      code[ 508] = 'h0000002300000000000000a500001500000000a40090160000000000008f2100;                                                                          // moveLong
      code[ 509] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 510] = 'h00000022000000000000000000a621000000008a000515000000000000000000;                                                                          // mov
      code[ 511] = 'h00000022000000000000000000a7210000000092000515000000000000000000;                                                                          // mov
      code[ 512] = 'h0000002300000000000000a700001500000000a60090160000000000008f2100;                                                                          // moveLong
      code[ 513] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 514] = 'h0000001f00000000000000000000010000000000003620000000000000000000;                                                                          // label
      code[ 515] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 516] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 517] = 'h0000002200000000000000920002150000000000009121000000000000000000;                                                                          // mov
      code[ 518] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 519] = 'h00000022000000000000000000a8210000000091000015000000000000000000;                                                                          // mov
      code[ 520] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 521] = 'h00000022000000000000008a0000150000000000008f21000000000000000000;                                                                          // mov
      code[ 522] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 523] = 'h00000022000000000000000000a9210000000091000615000000000000000000;                                                                          // mov
      code[ 524] = 'h00000022000000000000000000aa2100000000a900a816000000000000000000;                                                                          // mov
      code[ 525] = 'h0000001c000000000000001c003b21000000000000aa210000000000008a2100;                                                                          // jNe
      code[ 526] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 527] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 528] = 'h00000022000000000000000000ab21000000008a000515000000000000000000;                                                                          // mov
      code[ 529] = 'h00000022000000000000000000ac2100000000ab008f16000000000000000000;                                                                          // mov
      code[ 530] = 'h00000022000000000000000000ad210000000091000515000000000000000000;                                                                          // mov
      code[ 531] = 'h0000002200000000000000ad00a816000000000000ac21000000000000000000;                                                                          // mov
      code[ 532] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 533] = 'h00000022000000000000000000ae21000000008a000415000000000000000000;                                                                          // mov
      code[ 534] = 'h00000022000000000000000000af2100000000ae008f16000000000000000000;                                                                          // mov
      code[ 535] = 'h00000022000000000000000000b0210000000091000415000000000000000000;                                                                          // mov
      code[ 536] = 'h0000002200000000000000b000a816000000000000af21000000000000000000;                                                                          // mov
      code[ 537] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 538] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 539] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 540] = 'h00000022000000000000000000b121000000008a000415000000000000000000;                                                                          // mov
      code[ 541] = 'h00000030000000000000000000b1210000000000008f21000000000000062000;                                                                          // resize
      code[ 542] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 543] = 'h00000000000000000000000000b221000000000000a821000000000000012000;                                                                          // add
      code[ 544] = 'h000000220000000000000091000015000000000000b221000000000000000000;                                                                          // mov
      code[ 545] = 'h00000022000000000000000000b3210000000091000615000000000000000000;                                                                          // mov
      code[ 546] = 'h0000002200000000000000b300b2160000000000009221000000000000000000;                                                                          // mov
      code[ 547] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 548] = 'h00000022000000000000000000b421000000008a000515000000000000000000;                                                                          // mov
      code[ 549] = 'h00000030000000000000000000b4210000000000008f21000000000000072000;                                                                          // resize
      code[ 550] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 551] = 'h0000001e00000000000000d00031210000000000000000000000000000000000;                                                                          // jmp
      code[ 552] = 'h0000001e0000000000000026003c210000000000000000000000000000000000;                                                                          // jmp
      code[ 553] = 'h0000001f00000000000000000000010000000000003b20000000000000000000;                                                                          // label
      code[ 554] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 555] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 556] = 'h00000022000000000000000000b521000000008a000415000000000000000000;                                                                          // mov
      code[ 557] = 'h00000022000000000000000000b62100000000b5008f16000000000000000000;                                                                          // mov
      code[ 558] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 559] = 'h00000022000000000000000000b721000000008a000515000000000000000000;                                                                          // mov
      code[ 560] = 'h00000022000000000000000000b82100000000b7008f16000000000000000000;                                                                          // mov
      code[ 561] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 562] = 'h0000000e00000000000000000000010000000000009121000000000000002000;                                                                          // assertNe
      code[ 563] = 'h00000022000000000000000000b9210000000091000615000000000000000000;                                                                          // mov
      code[ 564] = 'h00000005000000000000000000ba21000000000000b9210000000000008a2100;                                                                          // arrayIndex
      code[ 565] = 'h00000038000000000000000000ba21000000000000ba21000000000000012000;                                                                          // subtract
      code[ 566] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 567] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 568] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 569] = 'h00000022000000000000000000bb21000000008a000515000000000000000000;                                                                          // mov
      code[ 570] = 'h00000030000000000000000000bb210000000000008f21000000000000072000;                                                                          // resize
      code[ 571] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 572] = 'h00000022000000000000000000bc21000000008a000415000000000000000000;                                                                          // mov
      code[ 573] = 'h00000030000000000000000000bc210000000000008f21000000000000062000;                                                                          // resize
      code[ 574] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 575] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 576] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 577] = 'h00000022000000000000000000bd210000000091000515000000000000000000;                                                                          // mov
      code[ 578] = 'h0000003700000000000000bd00ba16000000000000b821000000000000000000;                                                                          // shiftUp
      code[ 579] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 580] = 'h00000022000000000000000000be210000000091000415000000000000000000;                                                                          // mov
      code[ 581] = 'h0000003700000000000000be00ba16000000000000b621000000000000000000;                                                                          // shiftUp
      code[ 582] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 583] = 'h00000022000000000000000000bf210000000091000615000000000000000000;                                                                          // mov
      code[ 584] = 'h00000000000000000000000000c021000000000000ba21000000000000012000;                                                                          // add
      code[ 585] = 'h0000003700000000000000bf00c0160000000000009221000000000000000000;                                                                          // shiftUp
      code[ 586] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 587] = 'h0000000000000000000000910000150000000091000015000000000000012000;                                                                          // add
      code[ 588] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 589] = 'h0000001e00000000000000aa0031210000000000000000000000000000000000;                                                                          // jmp
      code[ 590] = 'h0000001f00000000000000000000010000000000003c20000000000000000000;                                                                          // label
      code[ 591] = 'h0000001f00000000000000000000010000000000003420000000000000000000;                                                                          // label
      code[ 592] = 'h00000001000000000000000000c1210000000000000520000000000000000000;                                                                          // array
      code[ 593] = 'h0000002200000000000000c10000150000000000008f21000000000000000000;                                                                          // mov
      code[ 594] = 'h0000002200000000000000c10002150000000000000020000000000000000000;                                                                          // mov
      code[ 595] = 'h00000001000000000000000000c2210000000000000620000000000000000000;                                                                          // array
      code[ 596] = 'h0000002200000000000000c1000415000000000000c221000000000000000000;                                                                          // mov
      code[ 597] = 'h00000001000000000000000000c3210000000000000720000000000000000000;                                                                          // array
      code[ 598] = 'h0000002200000000000000c1000515000000000000c321000000000000000000;                                                                          // mov
      code[ 599] = 'h0000002200000000000000c10006150000000000000020000000000000000000;                                                                          // mov
      code[ 600] = 'h0000002200000000000000c10003150000000000008d21000000000000000000;                                                                          // mov
      code[ 601] = 'h00000000000000000000008d000115000000008d000115000000000000012000;                                                                          // add
      code[ 602] = 'h0000002200000000000000c1000115000000008d000115000000000000000000;                                                                          // mov
      code[ 603] = 'h00000001000000000000000000c4210000000000000520000000000000000000;                                                                          // array
      code[ 604] = 'h0000002200000000000000c40000150000000000008f21000000000000000000;                                                                          // mov
      code[ 605] = 'h0000002200000000000000c40002150000000000000020000000000000000000;                                                                          // mov
      code[ 606] = 'h00000001000000000000000000c5210000000000000620000000000000000000;                                                                          // array
      code[ 607] = 'h0000002200000000000000c4000415000000000000c521000000000000000000;                                                                          // mov
      code[ 608] = 'h00000001000000000000000000c6210000000000000720000000000000000000;                                                                          // array
      code[ 609] = 'h0000002200000000000000c4000515000000000000c621000000000000000000;                                                                          // mov
      code[ 610] = 'h0000002200000000000000c40006150000000000000020000000000000000000;                                                                          // mov
      code[ 611] = 'h0000002200000000000000c40003150000000000008d21000000000000000000;                                                                          // mov
      code[ 612] = 'h00000000000000000000008d000115000000008d000115000000000000012000;                                                                          // add
      code[ 613] = 'h0000002200000000000000c4000115000000008d000115000000000000000000;                                                                          // mov
      code[ 614] = 'h00000025000000000000000000c721000000008a000615000000000000000000;                                                                          // not
      code[ 615] = 'h0000001c000000000000004c003d21000000000000c721000000000000002000;                                                                          // jNe
      code[ 616] = 'h00000001000000000000000000c8210000000000000820000000000000000000;                                                                          // array
      code[ 617] = 'h0000002200000000000000c1000615000000000000c821000000000000000000;                                                                          // mov
      code[ 618] = 'h00000001000000000000000000c9210000000000000820000000000000000000;                                                                          // array
      code[ 619] = 'h0000002200000000000000c4000615000000000000c921000000000000000000;                                                                          // mov
      code[ 620] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 621] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 622] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 623] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 624] = 'h00000022000000000000000000ca21000000008a000615000000000000000000;                                                                          // mov
      code[ 625] = 'h00000022000000000000000000cb2100000000c4000615000000000000000000;                                                                          // mov
      code[ 626] = 'h00000000000000000000000000cc210000000000008f21000000000000012000;                                                                          // add
      code[ 627] = 'h0000002300000000000000cb00001500000000ca009016000000000000cc2100;                                                                          // moveLong
      code[ 628] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 629] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 630] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 631] = 'h00000022000000000000000000cd21000000008a000515000000000000000000;                                                                          // mov
      code[ 632] = 'h00000022000000000000000000ce2100000000c4000515000000000000000000;                                                                          // mov
      code[ 633] = 'h0000002300000000000000ce00001500000000cd0090160000000000008f2100;                                                                          // moveLong
      code[ 634] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 635] = 'h00000022000000000000000000cf21000000008a000415000000000000000000;                                                                          // mov
      code[ 636] = 'h00000022000000000000000000d02100000000c4000415000000000000000000;                                                                          // mov
      code[ 637] = 'h0000002300000000000000d000001500000000cf0090160000000000008f2100;                                                                          // moveLong
      code[ 638] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 639] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 640] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 641] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 642] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 643] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 644] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 645] = 'h00000022000000000000000000d121000000008a000515000000000000000000;                                                                          // mov
      code[ 646] = 'h00000022000000000000000000d22100000000c1000515000000000000000000;                                                                          // mov
      code[ 647] = 'h0000002300000000000000d200001500000000d10000150000000000008f2100;                                                                          // moveLong
      code[ 648] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 649] = 'h00000022000000000000000000d321000000008a000415000000000000000000;                                                                          // mov
      code[ 650] = 'h00000022000000000000000000d42100000000c1000415000000000000000000;                                                                          // mov
      code[ 651] = 'h0000002300000000000000d400001500000000d30000150000000000008f2100;                                                                          // moveLong
      code[ 652] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 653] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 654] = 'h00000022000000000000000000d521000000008a000615000000000000000000;                                                                          // mov
      code[ 655] = 'h00000022000000000000000000d62100000000c1000615000000000000000000;                                                                          // mov
      code[ 656] = 'h00000000000000000000000000d7210000000000008f21000000000000012000;                                                                          // add
      code[ 657] = 'h0000002300000000000000d600001500000000d5000015000000000000d72100;                                                                          // moveLong
      code[ 658] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 659] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 660] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 661] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 662] = 'h00000022000000000000000000d82100000000c1000015000000000000000000;                                                                          // mov
      code[ 663] = 'h00000000000000000000000000d921000000000000d821000000000000012000;                                                                          // add
      code[ 664] = 'h00000022000000000000000000da2100000000c1000615000000000000000000;                                                                          // mov
      code[ 665] = 'h0000001f00000000000000000000010000000000003f20000000000000000000;                                                                          // label
      code[ 666] = 'h00000022000000000000000000db210000000000000020000000000000000000;                                                                          // mov
      code[ 667] = 'h0000001f00000000000000000000010000000000004020000000000000000000;                                                                          // label
      code[ 668] = 'h000000180000000000000006004221000000000000db21000000000000d92100;                                                                          // jGe
      code[ 669] = 'h00000022000000000000000000dc2100000000da00db16000000000000000000;                                                                          // mov
      code[ 670] = 'h0000002200000000000000dc000215000000000000c121000000000000000000;                                                                          // mov
      code[ 671] = 'h0000001f00000000000000000000010000000000004120000000000000000000;                                                                          // label
      code[ 672] = 'h00000000000000000000000000db21000000000000db21000000000000012000;                                                                          // add
      code[ 673] = 'h0000001e00000000fffffffa0040210000000000000000000000000000000000;                                                                          // jmp
      code[ 674] = 'h0000001f00000000000000000000010000000000004220000000000000000000;                                                                          // label
      code[ 675] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 676] = 'h00000022000000000000000000dd2100000000c4000015000000000000000000;                                                                          // mov
      code[ 677] = 'h00000000000000000000000000de21000000000000dd21000000000000012000;                                                                          // add
      code[ 678] = 'h00000022000000000000000000df2100000000c4000615000000000000000000;                                                                          // mov
      code[ 679] = 'h0000001f00000000000000000000010000000000004320000000000000000000;                                                                          // label
      code[ 680] = 'h00000022000000000000000000e0210000000000000020000000000000000000;                                                                          // mov
      code[ 681] = 'h0000001f00000000000000000000010000000000004420000000000000000000;                                                                          // label
      code[ 682] = 'h000000180000000000000006004621000000000000e021000000000000de2100;                                                                          // jGe
      code[ 683] = 'h00000022000000000000000000e12100000000df00e016000000000000000000;                                                                          // mov
      code[ 684] = 'h0000002200000000000000e1000215000000000000c421000000000000000000;                                                                          // mov
      code[ 685] = 'h0000001f00000000000000000000010000000000004520000000000000000000;                                                                          // label
      code[ 686] = 'h00000000000000000000000000e021000000000000e021000000000000012000;                                                                          // add
      code[ 687] = 'h0000001e00000000fffffffa0044210000000000000000000000000000000000;                                                                          // jmp
      code[ 688] = 'h0000001f00000000000000000000010000000000004620000000000000000000;                                                                          // label
      code[ 689] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 690] = 'h0000001e000000000000001d003e210000000000000000000000000000000000;                                                                          // jmp
      code[ 691] = 'h0000001f00000000000000000000010000000000003d20000000000000000000;                                                                          // label
      code[ 692] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 693] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 694] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 695] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 696] = 'h00000022000000000000000000e221000000008a000515000000000000000000;                                                                          // mov
      code[ 697] = 'h00000022000000000000000000e32100000000c1000515000000000000000000;                                                                          // mov
      code[ 698] = 'h0000002300000000000000e300001500000000e20000150000000000008f2100;                                                                          // moveLong
      code[ 699] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 700] = 'h00000022000000000000000000e421000000008a000415000000000000000000;                                                                          // mov
      code[ 701] = 'h00000022000000000000000000e52100000000c1000415000000000000000000;                                                                          // mov
      code[ 702] = 'h0000002300000000000000e500001500000000e40000150000000000008f2100;                                                                          // moveLong
      code[ 703] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 704] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 705] = 'h00000001000000000000000000e6210000000000000820000000000000000000;                                                                          // array
      code[ 706] = 'h00000022000000000000008a000615000000000000e621000000000000000000;                                                                          // mov
      code[ 707] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 708] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 709] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 710] = 'h00000022000000000000000000e721000000008a000515000000000000000000;                                                                          // mov
      code[ 711] = 'h00000022000000000000000000e82100000000c4000515000000000000000000;                                                                          // mov
      code[ 712] = 'h0000002300000000000000e800001500000000e70090160000000000008f2100;                                                                          // moveLong
      code[ 713] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 714] = 'h00000022000000000000000000e921000000008a000415000000000000000000;                                                                          // mov
      code[ 715] = 'h00000022000000000000000000ea2100000000c4000415000000000000000000;                                                                          // mov
      code[ 716] = 'h0000002300000000000000ea00001500000000e90090160000000000008f2100;                                                                          // moveLong
      code[ 717] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 718] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 719] = 'h0000001f00000000000000000000010000000000003e20000000000000000000;                                                                          // label
      code[ 720] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 721] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 722] = 'h0000002200000000000000c40002150000000000008a21000000000000000000;                                                                          // mov
      code[ 723] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 724] = 'h00000022000000000000000000eb21000000008a000415000000000000000000;                                                                          // mov
      code[ 725] = 'h00000022000000000000000000ec2100000000eb008f16000000000000000000;                                                                          // mov
      code[ 726] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 727] = 'h00000022000000000000000000ed21000000008a000515000000000000000000;                                                                          // mov
      code[ 728] = 'h00000022000000000000000000ee2100000000ed008f16000000000000000000;                                                                          // mov
      code[ 729] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 730] = 'h0000002200000000000000c10002150000000000008a21000000000000000000;                                                                          // mov
      code[ 731] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 732] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 733] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 734] = 'h00000022000000000000000000ef21000000008a000615000000000000000000;                                                                          // mov
      code[ 735] = 'h00000030000000000000000000ef210000000000000220000000000000082000;                                                                          // resize
      code[ 736] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 737] = 'h00000022000000000000000000f021000000008a000415000000000000000000;                                                                          // mov
      code[ 738] = 'h0000002200000000000000f0000015000000000000ec21000000000000000000;                                                                          // mov
      code[ 739] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 740] = 'h00000022000000000000008a0000150000000000000120000000000000000000;                                                                          // mov
      code[ 741] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 742] = 'h00000022000000000000000000f121000000008a000515000000000000000000;                                                                          // mov
      code[ 743] = 'h00000030000000000000000000f1210000000000000120000000000000072000;                                                                          // resize
      code[ 744] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 745] = 'h00000022000000000000000000f221000000008a000415000000000000000000;                                                                          // mov
      code[ 746] = 'h00000030000000000000000000f2210000000000000120000000000000062000;                                                                          // resize
      code[ 747] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 748] = 'h00000022000000000000000000f321000000008a000515000000000000000000;                                                                          // mov
      code[ 749] = 'h0000002200000000000000f3000015000000000000ee21000000000000000000;                                                                          // mov
      code[ 750] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 751] = 'h00000022000000000000000000f421000000008a000615000000000000000000;                                                                          // mov
      code[ 752] = 'h0000002200000000000000f4000015000000000000c121000000000000000000;                                                                          // mov
      code[ 753] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 754] = 'h00000022000000000000000000f521000000008a000615000000000000000000;                                                                          // mov
      code[ 755] = 'h0000002200000000000000f5000115000000000000c421000000000000000000;                                                                          // mov
      code[ 756] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 757] = 'h0000001e00000000000000020031210000000000000000000000000000000000;                                                                          // jmp
      code[ 758] = 'h0000001e00000000000000060033210000000000000000000000000000000000;                                                                          // jmp
      code[ 759] = 'h0000001f00000000000000000000010000000000003120000000000000000000;                                                                          // label
      code[ 760] = 'h000000220000000000000000008b210000000000000120000000000000000000;                                                                          // mov
      code[ 761] = 'h0000001e00000000000000030033210000000000000000000000000000000000;                                                                          // jmp
      code[ 762] = 'h0000001f00000000000000000000010000000000003220000000000000000000;                                                                          // label
      code[ 763] = 'h000000220000000000000000008b210000000000000020000000000000000000;                                                                          // mov
      code[ 764] = 'h0000001f00000000000000000000010000000000003320000000000000000000;                                                                          // label
      code[ 765] = 'h0000001c00000000000000020047210000000000008b21000000000000002000;                                                                          // jNe
      code[ 766] = 'h0000002200000000000000000017210000000000008a21000000000000000000;                                                                          // mov
      code[ 767] = 'h0000001f00000000000000000000010000000000004720000000000000000000;                                                                          // label
      code[ 768] = 'h0000001e0000000000000160002c210000000000000000000000000000000000;                                                                          // jmp
      code[ 769] = 'h0000001f00000000000000000000010000000000002e20000000000000000000;                                                                          // label
      code[ 770] = 'h00000022000000000000000000f6210000000017000415000000000000000000;                                                                          // mov
      code[ 771] = 'h00000005000000000000000000f721000000000000f621000000000000012100;                                                                          // arrayIndex
      code[ 772] = 'h000000160000000000000009004821000000000000f721000000000000002000;                                                                          // jEq
      code[ 773] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 774] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 775] = 'h0000002200000000000000030000150000000000001721000000000000000000;                                                                          // mov
      code[ 776] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 777] = 'h0000002200000000000000030001150000000000000120000000000000000000;                                                                          // mov
      code[ 778] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 779] = 'h000000380000000000000003000215000000000000f721000000000000012000;                                                                          // subtract
      code[ 780] = 'h0000001e000000000000015b0029210000000000000000000000000000000000;                                                                          // jmp
      code[ 781] = 'h0000001f00000000000000000000010000000000004820000000000000000000;                                                                          // label
      code[ 782] = 'h00000003000000000000000000f821000000000000f621000000000000012100;                                                                          // arrayCountLess
      code[ 783] = 'h00000025000000000000000000f9210000000017000615000000000000000000;                                                                          // not
      code[ 784] = 'h000000160000000000000009004921000000000000f921000000000000002000;                                                                          // jEq
      code[ 785] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 786] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 787] = 'h0000002200000000000000030000150000000000001721000000000000000000;                                                                          // mov
      code[ 788] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 789] = 'h0000002200000000000000030001150000000000000020000000000000000000;                                                                          // mov
      code[ 790] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 791] = 'h000000220000000000000003000215000000000000f821000000000000000000;                                                                          // mov
      code[ 792] = 'h0000001e000000000000014f0029210000000000000000000000000000000000;                                                                          // jmp
      code[ 793] = 'h0000001f00000000000000000000010000000000004920000000000000000000;                                                                          // label
      code[ 794] = 'h00000022000000000000000000fa210000000017000615000000000000000000;                                                                          // mov
      code[ 795] = 'h00000022000000000000000000fb2100000000fa00f816000000000000000000;                                                                          // mov
      code[ 796] = 'h0000001f00000000000000000000010000000000004a20000000000000000000;                                                                          // label
      code[ 797] = 'h00000022000000000000000000fd2100000000fb000015000000000000000000;                                                                          // mov
      code[ 798] = 'h00000022000000000000000000fe2100000000fb000315000000000000000000;                                                                          // mov
      code[ 799] = 'h00000022000000000000000000ff2100000000fe000215000000000000000000;                                                                          // mov
      code[ 800] = 'h0000001b000000000000013a004c21000000000000fd21000000000000ff2100;                                                                          // jLt
      code[ 801] = 'h000000220000000000000000010021000000000000ff21000000000000000000;                                                                          // mov
      code[ 802] = 'h0000003600000000000000000100210000000000000120000000000000000000;                                                                          // shiftRight
      code[ 803] = 'h0000000000000000000000000101210000000000010021000000000000012000;                                                                          // add
      code[ 804] = 'h00000022000000000000000001022100000000fb000215000000000000000000;                                                                          // mov
      code[ 805] = 'h00000016000000000000008a004e210000000000010221000000000000002000;                                                                          // jEq
      code[ 806] = 'h0000000100000000000000000103210000000000000520000000000000000000;                                                                          // array
      code[ 807] = 'h0000002200000000000001030000150000000000010021000000000000000000;                                                                          // mov
      code[ 808] = 'h0000002200000000000001030002150000000000000020000000000000000000;                                                                          // mov
      code[ 809] = 'h0000000100000000000000000104210000000000000620000000000000000000;                                                                          // array
      code[ 810] = 'h0000002200000000000001030004150000000000010421000000000000000000;                                                                          // mov
      code[ 811] = 'h0000000100000000000000000105210000000000000720000000000000000000;                                                                          // array
      code[ 812] = 'h0000002200000000000001030005150000000000010521000000000000000000;                                                                          // mov
      code[ 813] = 'h0000002200000000000001030006150000000000000020000000000000000000;                                                                          // mov
      code[ 814] = 'h000000220000000000000103000315000000000000fe21000000000000000000;                                                                          // mov
      code[ 815] = 'h0000000000000000000000fe00011500000000fe000115000000000000012000;                                                                          // add
      code[ 816] = 'h00000022000000000000010300011500000000fe000115000000000000000000;                                                                          // mov
      code[ 817] = 'h00000025000000000000000001062100000000fb000615000000000000000000;                                                                          // not
      code[ 818] = 'h0000001c0000000000000025004f210000000000010621000000000000002000;                                                                          // jNe
      code[ 819] = 'h0000000100000000000000000107210000000000000820000000000000000000;                                                                          // array
      code[ 820] = 'h0000002200000000000001030006150000000000010721000000000000000000;                                                                          // mov
      code[ 821] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 822] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 823] = 'h00000022000000000000000001082100000000fb000615000000000000000000;                                                                          // mov
      code[ 824] = 'h0000002200000000000000000109210000000103000615000000000000000000;                                                                          // mov
      code[ 825] = 'h000000000000000000000000010a210000000000010021000000000000012000;                                                                          // add
      code[ 826] = 'h00000023000000000000010900001500000001080101160000000000010a2100;                                                                          // moveLong
      code[ 827] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 828] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 829] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 830] = 'h000000220000000000000000010b2100000000fb000415000000000000000000;                                                                          // mov
      code[ 831] = 'h000000220000000000000000010c210000000103000415000000000000000000;                                                                          // mov
      code[ 832] = 'h00000023000000000000010c000015000000010b010116000000000001002100;                                                                          // moveLong
      code[ 833] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 834] = 'h000000220000000000000000010d2100000000fb000515000000000000000000;                                                                          // mov
      code[ 835] = 'h000000220000000000000000010e210000000103000515000000000000000000;                                                                          // mov
      code[ 836] = 'h00000023000000000000010e000015000000010d010116000000000001002100;                                                                          // moveLong
      code[ 837] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 838] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 839] = 'h000000220000000000000000010f210000000103000015000000000000000000;                                                                          // mov
      code[ 840] = 'h0000000000000000000000000110210000000000010f21000000000000012000;                                                                          // add
      code[ 841] = 'h0000002200000000000000000111210000000103000615000000000000000000;                                                                          // mov
      code[ 842] = 'h0000001f00000000000000000000010000000000005120000000000000000000;                                                                          // label
      code[ 843] = 'h0000002200000000000000000112210000000000000020000000000000000000;                                                                          // mov
      code[ 844] = 'h0000001f00000000000000000000010000000000005220000000000000000000;                                                                          // label
      code[ 845] = 'h0000001800000000000000060054210000000000011221000000000001102100;                                                                          // jGe
      code[ 846] = 'h0000002200000000000000000113210000000111011216000000000000000000;                                                                          // mov
      code[ 847] = 'h0000002200000000000001130002150000000000010321000000000000000000;                                                                          // mov
      code[ 848] = 'h0000001f00000000000000000000010000000000005320000000000000000000;                                                                          // label
      code[ 849] = 'h0000000000000000000000000112210000000000011221000000000000012000;                                                                          // add
      code[ 850] = 'h0000001e00000000fffffffa0052210000000000000000000000000000000000;                                                                          // jmp
      code[ 851] = 'h0000001f00000000000000000000010000000000005420000000000000000000;                                                                          // label
      code[ 852] = 'h00000022000000000000000001142100000000fb000615000000000000000000;                                                                          // mov
      code[ 853] = 'h0000003000000000000000000114210000000000010121000000000000082000;                                                                          // resize
      code[ 854] = 'h0000001e000000000000000c0050210000000000000000000000000000000000;                                                                          // jmp
      code[ 855] = 'h0000001f00000000000000000000010000000000004f20000000000000000000;                                                                          // label
      code[ 856] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 857] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 858] = 'h00000022000000000000000001152100000000fb000415000000000000000000;                                                                          // mov
      code[ 859] = 'h0000002200000000000000000116210000000103000415000000000000000000;                                                                          // mov
      code[ 860] = 'h0000002300000000000001160000150000000115010116000000000001002100;                                                                          // moveLong
      code[ 861] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 862] = 'h00000022000000000000000001172100000000fb000515000000000000000000;                                                                          // mov
      code[ 863] = 'h0000002200000000000000000118210000000103000515000000000000000000;                                                                          // mov
      code[ 864] = 'h0000002300000000000001180000150000000117010116000000000001002100;                                                                          // moveLong
      code[ 865] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 866] = 'h0000001f00000000000000000000010000000000005020000000000000000000;                                                                          // label
      code[ 867] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 868] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 869] = 'h0000002200000000000001030002150000000000010221000000000000000000;                                                                          // mov
      code[ 870] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 871] = 'h0000002200000000000000000119210000000102000015000000000000000000;                                                                          // mov
      code[ 872] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 873] = 'h0000002200000000000000fb0000150000000000010021000000000000000000;                                                                          // mov
      code[ 874] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 875] = 'h000000220000000000000000011a210000000102000615000000000000000000;                                                                          // mov
      code[ 876] = 'h000000220000000000000000011b21000000011a011916000000000000000000;                                                                          // mov
      code[ 877] = 'h0000001c000000000000001c0055210000000000011b21000000000000fb2100;                                                                          // jNe
      code[ 878] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 879] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 880] = 'h000000220000000000000000011c2100000000fb000515000000000000000000;                                                                          // mov
      code[ 881] = 'h000000220000000000000000011d21000000011c010016000000000000000000;                                                                          // mov
      code[ 882] = 'h000000220000000000000000011e210000000102000515000000000000000000;                                                                          // mov
      code[ 883] = 'h00000022000000000000011e0119160000000000011d21000000000000000000;                                                                          // mov
      code[ 884] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 885] = 'h000000220000000000000000011f2100000000fb000415000000000000000000;                                                                          // mov
      code[ 886] = 'h000000220000000000000000012021000000011f010016000000000000000000;                                                                          // mov
      code[ 887] = 'h0000002200000000000000000121210000000102000415000000000000000000;                                                                          // mov
      code[ 888] = 'h0000002200000000000001210119160000000000012021000000000000000000;                                                                          // mov
      code[ 889] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 890] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 891] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 892] = 'h00000022000000000000000001222100000000fb000515000000000000000000;                                                                          // mov
      code[ 893] = 'h0000003000000000000000000122210000000000010021000000000000072000;                                                                          // resize
      code[ 894] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 895] = 'h00000022000000000000000001232100000000fb000415000000000000000000;                                                                          // mov
      code[ 896] = 'h0000003000000000000000000123210000000000010021000000000000062000;                                                                          // resize
      code[ 897] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 898] = 'h0000000000000000000000000124210000000000011921000000000000012000;                                                                          // add
      code[ 899] = 'h0000002200000000000001020000150000000000012421000000000000000000;                                                                          // mov
      code[ 900] = 'h0000002200000000000000000125210000000102000615000000000000000000;                                                                          // mov
      code[ 901] = 'h0000002200000000000001250124160000000000010321000000000000000000;                                                                          // mov
      code[ 902] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 903] = 'h0000001e00000000000000d0004b210000000000000000000000000000000000;                                                                          // jmp
      code[ 904] = 'h0000001e00000000000000260056210000000000000000000000000000000000;                                                                          // jmp
      code[ 905] = 'h0000001f00000000000000000000010000000000005520000000000000000000;                                                                          // label
      code[ 906] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 907] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 908] = 'h0000000e00000000000000000000010000000000010221000000000000002000;                                                                          // assertNe
      code[ 909] = 'h0000002200000000000000000126210000000102000615000000000000000000;                                                                          // mov
      code[ 910] = 'h0000000500000000000000000127210000000000012621000000000000fb2100;                                                                          // arrayIndex
      code[ 911] = 'h0000003800000000000000000127210000000000012721000000000000012000;                                                                          // subtract
      code[ 912] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 913] = 'h00000022000000000000000001282100000000fb000515000000000000000000;                                                                          // mov
      code[ 914] = 'h0000002200000000000000000129210000000128010016000000000000000000;                                                                          // mov
      code[ 915] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 916] = 'h000000220000000000000000012a2100000000fb000415000000000000000000;                                                                          // mov
      code[ 917] = 'h000000220000000000000000012b21000000012a010016000000000000000000;                                                                          // mov
      code[ 918] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 919] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 920] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 921] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 922] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 923] = 'h000000220000000000000000012c210000000102000515000000000000000000;                                                                          // mov
      code[ 924] = 'h00000037000000000000012c0127160000000000012921000000000000000000;                                                                          // shiftUp
      code[ 925] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 926] = 'h000000220000000000000000012d210000000102000615000000000000000000;                                                                          // mov
      code[ 927] = 'h000000000000000000000000012e210000000000012721000000000000012000;                                                                          // add
      code[ 928] = 'h00000037000000000000012d012e160000000000010321000000000000000000;                                                                          // shiftUp
      code[ 929] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 930] = 'h000000220000000000000000012f210000000102000415000000000000000000;                                                                          // mov
      code[ 931] = 'h00000037000000000000012f0127160000000000012b21000000000000000000;                                                                          // shiftUp
      code[ 932] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 933] = 'h0000000000000000000001020000150000000102000015000000000000012000;                                                                          // add
      code[ 934] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 935] = 'h00000022000000000000000001302100000000fb000415000000000000000000;                                                                          // mov
      code[ 936] = 'h0000003000000000000000000130210000000000010021000000000000062000;                                                                          // resize
      code[ 937] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 938] = 'h00000022000000000000000001312100000000fb000515000000000000000000;                                                                          // mov
      code[ 939] = 'h0000003000000000000000000131210000000000010021000000000000072000;                                                                          // resize
      code[ 940] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 941] = 'h0000001e00000000000000aa004b210000000000000000000000000000000000;                                                                          // jmp
      code[ 942] = 'h0000001f00000000000000000000010000000000005620000000000000000000;                                                                          // label
      code[ 943] = 'h0000001f00000000000000000000010000000000004e20000000000000000000;                                                                          // label
      code[ 944] = 'h0000000100000000000000000132210000000000000520000000000000000000;                                                                          // array
      code[ 945] = 'h0000002200000000000001320000150000000000010021000000000000000000;                                                                          // mov
      code[ 946] = 'h0000002200000000000001320002150000000000000020000000000000000000;                                                                          // mov
      code[ 947] = 'h0000000100000000000000000133210000000000000620000000000000000000;                                                                          // array
      code[ 948] = 'h0000002200000000000001320004150000000000013321000000000000000000;                                                                          // mov
      code[ 949] = 'h0000000100000000000000000134210000000000000720000000000000000000;                                                                          // array
      code[ 950] = 'h0000002200000000000001320005150000000000013421000000000000000000;                                                                          // mov
      code[ 951] = 'h0000002200000000000001320006150000000000000020000000000000000000;                                                                          // mov
      code[ 952] = 'h000000220000000000000132000315000000000000fe21000000000000000000;                                                                          // mov
      code[ 953] = 'h0000000000000000000000fe00011500000000fe000115000000000000012000;                                                                          // add
      code[ 954] = 'h00000022000000000000013200011500000000fe000115000000000000000000;                                                                          // mov
      code[ 955] = 'h0000000100000000000000000135210000000000000520000000000000000000;                                                                          // array
      code[ 956] = 'h0000002200000000000001350000150000000000010021000000000000000000;                                                                          // mov
      code[ 957] = 'h0000002200000000000001350002150000000000000020000000000000000000;                                                                          // mov
      code[ 958] = 'h0000000100000000000000000136210000000000000620000000000000000000;                                                                          // array
      code[ 959] = 'h0000002200000000000001350004150000000000013621000000000000000000;                                                                          // mov
      code[ 960] = 'h0000000100000000000000000137210000000000000720000000000000000000;                                                                          // array
      code[ 961] = 'h0000002200000000000001350005150000000000013721000000000000000000;                                                                          // mov
      code[ 962] = 'h0000002200000000000001350006150000000000000020000000000000000000;                                                                          // mov
      code[ 963] = 'h000000220000000000000135000315000000000000fe21000000000000000000;                                                                          // mov
      code[ 964] = 'h0000000000000000000000fe00011500000000fe000115000000000000012000;                                                                          // add
      code[ 965] = 'h00000022000000000000013500011500000000fe000115000000000000000000;                                                                          // mov
      code[ 966] = 'h00000025000000000000000001382100000000fb000615000000000000000000;                                                                          // not
      code[ 967] = 'h0000001c000000000000004c0057210000000000013821000000000000002000;                                                                          // jNe
      code[ 968] = 'h0000000100000000000000000139210000000000000820000000000000000000;                                                                          // array
      code[ 969] = 'h0000002200000000000001320006150000000000013921000000000000000000;                                                                          // mov
      code[ 970] = 'h000000010000000000000000013a210000000000000820000000000000000000;                                                                          // array
      code[ 971] = 'h0000002200000000000001350006150000000000013a21000000000000000000;                                                                          // mov
      code[ 972] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 973] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 974] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 975] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 976] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 977] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 978] = 'h000000220000000000000000013b2100000000fb000515000000000000000000;                                                                          // mov
      code[ 979] = 'h000000220000000000000000013c210000000132000515000000000000000000;                                                                          // mov
      code[ 980] = 'h00000023000000000000013c000015000000013b000015000000000001002100;                                                                          // moveLong
      code[ 981] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 982] = 'h000000220000000000000000013d2100000000fb000415000000000000000000;                                                                          // mov
      code[ 983] = 'h000000220000000000000000013e210000000132000415000000000000000000;                                                                          // mov
      code[ 984] = 'h00000023000000000000013e000015000000013d000015000000000001002100;                                                                          // moveLong
      code[ 985] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 986] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 987] = 'h000000220000000000000000013f2100000000fb000615000000000000000000;                                                                          // mov
      code[ 988] = 'h0000002200000000000000000140210000000132000615000000000000000000;                                                                          // mov
      code[ 989] = 'h0000000000000000000000000141210000000000010021000000000000012000;                                                                          // add
      code[ 990] = 'h000000230000000000000140000015000000013f000015000000000001412100;                                                                          // moveLong
      code[ 991] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[ 992] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 993] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[ 994] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[ 995] = 'h00000022000000000000000001422100000000fb000615000000000000000000;                                                                          // mov
      code[ 996] = 'h0000002200000000000000000143210000000135000615000000000000000000;                                                                          // mov
      code[ 997] = 'h0000000000000000000000000144210000000000010021000000000000012000;                                                                          // add
      code[ 998] = 'h0000002300000000000001430000150000000142010116000000000001442100;                                                                          // moveLong
      code[ 999] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1000] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1001] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1002] = 'h00000022000000000000000001452100000000fb000515000000000000000000;                                                                          // mov
      code[1003] = 'h0000002200000000000000000146210000000135000515000000000000000000;                                                                          // mov
      code[1004] = 'h0000002300000000000001460000150000000145010116000000000001002100;                                                                          // moveLong
      code[1005] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1006] = 'h00000022000000000000000001472100000000fb000415000000000000000000;                                                                          // mov
      code[1007] = 'h0000002200000000000000000148210000000135000415000000000000000000;                                                                          // mov
      code[1008] = 'h0000002300000000000001480000150000000147010116000000000001002100;                                                                          // moveLong
      code[1009] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1010] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1011] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1012] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1013] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1014] = 'h0000002200000000000000000149210000000132000015000000000000000000;                                                                          // mov
      code[1015] = 'h000000000000000000000000014a210000000000014921000000000000012000;                                                                          // add
      code[1016] = 'h000000220000000000000000014b210000000132000615000000000000000000;                                                                          // mov
      code[1017] = 'h0000001f00000000000000000000010000000000005920000000000000000000;                                                                          // label
      code[1018] = 'h000000220000000000000000014c210000000000000020000000000000000000;                                                                          // mov
      code[1019] = 'h0000001f00000000000000000000010000000000005a20000000000000000000;                                                                          // label
      code[1020] = 'h000000180000000000000006005c210000000000014c210000000000014a2100;                                                                          // jGe
      code[1021] = 'h000000220000000000000000014d21000000014b014c16000000000000000000;                                                                          // mov
      code[1022] = 'h00000022000000000000014d0002150000000000013221000000000000000000;                                                                          // mov
      code[1023] = 'h0000001f00000000000000000000010000000000005b20000000000000000000;                                                                          // label
      code[1024] = 'h000000000000000000000000014c210000000000014c21000000000000012000;                                                                          // add
      code[1025] = 'h0000001e00000000fffffffa005a210000000000000000000000000000000000;                                                                          // jmp
      code[1026] = 'h0000001f00000000000000000000010000000000005c20000000000000000000;                                                                          // label
      code[1027] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1028] = 'h000000220000000000000000014e210000000135000015000000000000000000;                                                                          // mov
      code[1029] = 'h000000000000000000000000014f210000000000014e21000000000000012000;                                                                          // add
      code[1030] = 'h0000002200000000000000000150210000000135000615000000000000000000;                                                                          // mov
      code[1031] = 'h0000001f00000000000000000000010000000000005d20000000000000000000;                                                                          // label
      code[1032] = 'h0000002200000000000000000151210000000000000020000000000000000000;                                                                          // mov
      code[1033] = 'h0000001f00000000000000000000010000000000005e20000000000000000000;                                                                          // label
      code[1034] = 'h00000018000000000000000600602100000000000151210000000000014f2100;                                                                          // jGe
      code[1035] = 'h0000002200000000000000000152210000000150015116000000000000000000;                                                                          // mov
      code[1036] = 'h0000002200000000000001520002150000000000013521000000000000000000;                                                                          // mov
      code[1037] = 'h0000001f00000000000000000000010000000000005f20000000000000000000;                                                                          // label
      code[1038] = 'h0000000000000000000000000151210000000000015121000000000000012000;                                                                          // add
      code[1039] = 'h0000001e00000000fffffffa005e210000000000000000000000000000000000;                                                                          // jmp
      code[1040] = 'h0000001f00000000000000000000010000000000006020000000000000000000;                                                                          // label
      code[1041] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1042] = 'h0000001e000000000000001d0058210000000000000000000000000000000000;                                                                          // jmp
      code[1043] = 'h0000001f00000000000000000000010000000000005720000000000000000000;                                                                          // label
      code[1044] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1045] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1046] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1047] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1048] = 'h00000022000000000000000001532100000000fb000515000000000000000000;                                                                          // mov
      code[1049] = 'h0000002200000000000000000154210000000135000515000000000000000000;                                                                          // mov
      code[1050] = 'h0000002300000000000001540000150000000153010116000000000001002100;                                                                          // moveLong
      code[1051] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1052] = 'h00000022000000000000000001552100000000fb000415000000000000000000;                                                                          // mov
      code[1053] = 'h0000002200000000000000000156210000000135000415000000000000000000;                                                                          // mov
      code[1054] = 'h0000002300000000000001560000150000000155010116000000000001002100;                                                                          // moveLong
      code[1055] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1056] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1057] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1058] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1059] = 'h00000022000000000000000001572100000000fb000415000000000000000000;                                                                          // mov
      code[1060] = 'h0000002200000000000000000158210000000132000415000000000000000000;                                                                          // mov
      code[1061] = 'h0000002300000000000001580000150000000157000015000000000001002100;                                                                          // moveLong
      code[1062] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1063] = 'h00000022000000000000000001592100000000fb000515000000000000000000;                                                                          // mov
      code[1064] = 'h000000220000000000000000015a210000000132000515000000000000000000;                                                                          // mov
      code[1065] = 'h00000023000000000000015a0000150000000159000015000000000001002100;                                                                          // moveLong
      code[1066] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1067] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1068] = 'h000000010000000000000000015b210000000000000820000000000000000000;                                                                          // array
      code[1069] = 'h0000002200000000000000fb0006150000000000015b21000000000000000000;                                                                          // mov
      code[1070] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1071] = 'h0000001f00000000000000000000010000000000005820000000000000000000;                                                                          // label
      code[1072] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1073] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1074] = 'h000000220000000000000135000215000000000000fb21000000000000000000;                                                                          // mov
      code[1075] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1076] = 'h000000220000000000000000015c2100000000fb000415000000000000000000;                                                                          // mov
      code[1077] = 'h000000220000000000000000015d21000000015c010016000000000000000000;                                                                          // mov
      code[1078] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1079] = 'h000000220000000000000000015e2100000000fb000515000000000000000000;                                                                          // mov
      code[1080] = 'h000000220000000000000000015f21000000015e010016000000000000000000;                                                                          // mov
      code[1081] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1082] = 'h000000220000000000000132000215000000000000fb21000000000000000000;                                                                          // mov
      code[1083] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1084] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1085] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1086] = 'h00000022000000000000000001602100000000fb000615000000000000000000;                                                                          // mov
      code[1087] = 'h0000002200000000000001600000150000000000013221000000000000000000;                                                                          // mov
      code[1088] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1089] = 'h00000022000000000000000001612100000000fb000515000000000000000000;                                                                          // mov
      code[1090] = 'h0000002200000000000001610000150000000000015f21000000000000000000;                                                                          // mov
      code[1091] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1092] = 'h00000022000000000000000001622100000000fb000415000000000000000000;                                                                          // mov
      code[1093] = 'h0000002200000000000001620000150000000000015d21000000000000000000;                                                                          // mov
      code[1094] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1095] = 'h00000022000000000000000001632100000000fb000415000000000000000000;                                                                          // mov
      code[1096] = 'h0000003000000000000000000163210000000000000120000000000000062000;                                                                          // resize
      code[1097] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1098] = 'h00000022000000000000000001642100000000fb000615000000000000000000;                                                                          // mov
      code[1099] = 'h0000002200000000000001640001150000000000013521000000000000000000;                                                                          // mov
      code[1100] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1101] = 'h00000022000000000000000001652100000000fb000515000000000000000000;                                                                          // mov
      code[1102] = 'h0000003000000000000000000165210000000000000120000000000000072000;                                                                          // resize
      code[1103] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1104] = 'h0000002200000000000000fb0000150000000000000120000000000000000000;                                                                          // mov
      code[1105] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1106] = 'h00000022000000000000000001662100000000fb000615000000000000000000;                                                                          // mov
      code[1107] = 'h0000003000000000000000000166210000000000000220000000000000082000;                                                                          // resize
      code[1108] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1109] = 'h0000001e0000000000000002004b210000000000000000000000000000000000;                                                                          // jmp
      code[1110] = 'h0000001e0000000000000006004d210000000000000000000000000000000000;                                                                          // jmp
      code[1111] = 'h0000001f00000000000000000000010000000000004b20000000000000000000;                                                                          // label
      code[1112] = 'h00000022000000000000000000fc210000000000000120000000000000000000;                                                                          // mov
      code[1113] = 'h0000001e0000000000000003004d210000000000000000000000000000000000;                                                                          // jmp
      code[1114] = 'h0000001f00000000000000000000010000000000004c20000000000000000000;                                                                          // label
      code[1115] = 'h00000022000000000000000000fc210000000000000020000000000000000000;                                                                          // mov
      code[1116] = 'h0000001f00000000000000000000010000000000004d20000000000000000000;                                                                          // label
      code[1117] = 'h0000001c0000000000000002006121000000000000fc21000000000000002000;                                                                          // jNe
      code[1118] = 'h000000220000000000000000001721000000000000fb21000000000000000000;                                                                          // mov
      code[1119] = 'h0000001f00000000000000000000010000000000006120000000000000000000;                                                                          // label
      code[1120] = 'h0000001f00000000000000000000010000000000002c20000000000000000000;                                                                          // label
      code[1121] = 'h0000000000000000000000000083210000000000008321000000000000012000;                                                                          // add
      code[1122] = 'h0000001e00000000fffffd46002b210000000000000000000000000000000000;                                                                          // jmp
      code[1123] = 'h0000001f00000000000000000000010000000000002d20000000000000000000;                                                                          // label
      code[1124] = 'h0000000700000000000000000000010000000000000000000000000000000000;                                                                          // assert
      code[1125] = 'h0000001f00000000000000000000010000000000002720000000000000000000;                                                                          // label
      code[1126] = 'h0000001f00000000000000000000010000000000002820000000000000000000;                                                                          // label
      code[1127] = 'h0000001f00000000000000000000010000000000002920000000000000000000;                                                                          // label
      code[1128] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1129] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1130] = 'h0000002200000000000000000167210000000003000015000000000000000000;                                                                          // mov
      code[1131] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1132] = 'h0000002200000000000000000168210000000003000115000000000000000000;                                                                          // mov
      code[1133] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1134] = 'h0000002200000000000000000169210000000003000215000000000000000000;                                                                          // mov
      code[1135] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1136] = 'h0000001c00000000000000040062210000000000016821000000000000012000;                                                                          // jNe
      code[1137] = 'h000000220000000000000000016a210000000167000515000000000000000000;                                                                          // mov
      code[1138] = 'h00000022000000000000016a0169160000000000000121000000000000000000;                                                                          // mov
      code[1139] = 'h0000001e000000000000015d0008210000000000000000000000000000000000;                                                                          // jmp
      code[1140] = 'h0000001f00000000000000000000010000000000006220000000000000000000;                                                                          // label
      code[1141] = 'h0000001c000000000000000c0063210000000000016821000000000000022000;                                                                          // jNe
      code[1142] = 'h000000000000000000000000016b210000000000016921000000000000012000;                                                                          // add
      code[1143] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1144] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1145] = 'h000000220000000000000000016c210000000167000515000000000000000000;                                                                          // mov
      code[1146] = 'h00000037000000000000016c016b160000000000000121000000000000000000;                                                                          // shiftUp
      code[1147] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1148] = 'h000000220000000000000000016d210000000167000415000000000000000000;                                                                          // mov
      code[1149] = 'h00000037000000000000016d016b160000000000000121000000000000000000;                                                                          // shiftUp
      code[1150] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1151] = 'h0000000000000000000001670000150000000167000015000000000000012000;                                                                          // add
      code[1152] = 'h0000001e000000000000000b0064210000000000000000000000000000000000;                                                                          // jmp
      code[1153] = 'h0000001f00000000000000000000010000000000006320000000000000000000;                                                                          // label
      code[1154] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1155] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1156] = 'h000000220000000000000000016e210000000167000415000000000000000000;                                                                          // mov
      code[1157] = 'h00000037000000000000016e0169160000000000000121000000000000000000;                                                                          // shiftUp
      code[1158] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1159] = 'h000000220000000000000000016f210000000167000515000000000000000000;                                                                          // mov
      code[1160] = 'h00000037000000000000016f0169160000000000000121000000000000000000;                                                                          // shiftUp
      code[1161] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1162] = 'h0000000000000000000001670000150000000167000015000000000000012000;                                                                          // add
      code[1163] = 'h0000001f00000000000000000000010000000000006420000000000000000000;                                                                          // label
      code[1164] = 'h0000000000000000000000000000150000000000000015000000000000012000;                                                                          // add
      code[1165] = 'h0000001f00000000000000000000010000000000006520000000000000000000;                                                                          // label
      code[1166] = 'h0000002200000000000000000171210000000167000015000000000000000000;                                                                          // mov
      code[1167] = 'h0000002200000000000000000172210000000167000315000000000000000000;                                                                          // mov
      code[1168] = 'h0000002200000000000000000173210000000172000215000000000000000000;                                                                          // mov
      code[1169] = 'h0000001b000000000000013a0067210000000000017121000000000001732100;                                                                          // jLt
      code[1170] = 'h0000002200000000000000000174210000000000017321000000000000000000;                                                                          // mov
      code[1171] = 'h0000003600000000000000000174210000000000000120000000000000000000;                                                                          // shiftRight
      code[1172] = 'h0000000000000000000000000175210000000000017421000000000000012000;                                                                          // add
      code[1173] = 'h0000002200000000000000000176210000000167000215000000000000000000;                                                                          // mov
      code[1174] = 'h00000016000000000000008a0069210000000000017621000000000000002000;                                                                          // jEq
      code[1175] = 'h0000000100000000000000000177210000000000000520000000000000000000;                                                                          // array
      code[1176] = 'h0000002200000000000001770000150000000000017421000000000000000000;                                                                          // mov
      code[1177] = 'h0000002200000000000001770002150000000000000020000000000000000000;                                                                          // mov
      code[1178] = 'h0000000100000000000000000178210000000000000620000000000000000000;                                                                          // array
      code[1179] = 'h0000002200000000000001770004150000000000017821000000000000000000;                                                                          // mov
      code[1180] = 'h0000000100000000000000000179210000000000000720000000000000000000;                                                                          // array
      code[1181] = 'h0000002200000000000001770005150000000000017921000000000000000000;                                                                          // mov
      code[1182] = 'h0000002200000000000001770006150000000000000020000000000000000000;                                                                          // mov
      code[1183] = 'h0000002200000000000001770003150000000000017221000000000000000000;                                                                          // mov
      code[1184] = 'h0000000000000000000001720001150000000172000115000000000000012000;                                                                          // add
      code[1185] = 'h0000002200000000000001770001150000000172000115000000000000000000;                                                                          // mov
      code[1186] = 'h000000250000000000000000017a210000000167000615000000000000000000;                                                                          // not
      code[1187] = 'h0000001c0000000000000025006a210000000000017a21000000000000002000;                                                                          // jNe
      code[1188] = 'h000000010000000000000000017b210000000000000820000000000000000000;                                                                          // array
      code[1189] = 'h0000002200000000000001770006150000000000017b21000000000000000000;                                                                          // mov
      code[1190] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1191] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1192] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1193] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1194] = 'h000000220000000000000000017c210000000167000515000000000000000000;                                                                          // mov
      code[1195] = 'h000000220000000000000000017d210000000177000515000000000000000000;                                                                          // mov
      code[1196] = 'h00000023000000000000017d000015000000017c017516000000000001742100;                                                                          // moveLong
      code[1197] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1198] = 'h000000220000000000000000017e210000000167000415000000000000000000;                                                                          // mov
      code[1199] = 'h000000220000000000000000017f210000000177000415000000000000000000;                                                                          // mov
      code[1200] = 'h00000023000000000000017f000015000000017e017516000000000001742100;                                                                          // moveLong
      code[1201] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1202] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1203] = 'h0000002200000000000000000180210000000167000615000000000000000000;                                                                          // mov
      code[1204] = 'h0000002200000000000000000181210000000177000615000000000000000000;                                                                          // mov
      code[1205] = 'h0000000000000000000000000182210000000000017421000000000000012000;                                                                          // add
      code[1206] = 'h0000002300000000000001810000150000000180017516000000000001822100;                                                                          // moveLong
      code[1207] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1208] = 'h0000002200000000000000000183210000000177000015000000000000000000;                                                                          // mov
      code[1209] = 'h0000000000000000000000000184210000000000018321000000000000012000;                                                                          // add
      code[1210] = 'h0000002200000000000000000185210000000177000615000000000000000000;                                                                          // mov
      code[1211] = 'h0000001f00000000000000000000010000000000006c20000000000000000000;                                                                          // label
      code[1212] = 'h0000002200000000000000000186210000000000000020000000000000000000;                                                                          // mov
      code[1213] = 'h0000001f00000000000000000000010000000000006d20000000000000000000;                                                                          // label
      code[1214] = 'h000000180000000000000006006f210000000000018621000000000001842100;                                                                          // jGe
      code[1215] = 'h0000002200000000000000000187210000000185018616000000000000000000;                                                                          // mov
      code[1216] = 'h0000002200000000000001870002150000000000017721000000000000000000;                                                                          // mov
      code[1217] = 'h0000001f00000000000000000000010000000000006e20000000000000000000;                                                                          // label
      code[1218] = 'h0000000000000000000000000186210000000000018621000000000000012000;                                                                          // add
      code[1219] = 'h0000001e00000000fffffffa006d210000000000000000000000000000000000;                                                                          // jmp
      code[1220] = 'h0000001f00000000000000000000010000000000006f20000000000000000000;                                                                          // label
      code[1221] = 'h0000002200000000000000000188210000000167000615000000000000000000;                                                                          // mov
      code[1222] = 'h0000003000000000000000000188210000000000017521000000000000082000;                                                                          // resize
      code[1223] = 'h0000001e000000000000000c006b210000000000000000000000000000000000;                                                                          // jmp
      code[1224] = 'h0000001f00000000000000000000010000000000006a20000000000000000000;                                                                          // label
      code[1225] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1226] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1227] = 'h0000002200000000000000000189210000000167000415000000000000000000;                                                                          // mov
      code[1228] = 'h000000220000000000000000018a210000000177000415000000000000000000;                                                                          // mov
      code[1229] = 'h00000023000000000000018a0000150000000189017516000000000001742100;                                                                          // moveLong
      code[1230] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1231] = 'h000000220000000000000000018b210000000167000515000000000000000000;                                                                          // mov
      code[1232] = 'h000000220000000000000000018c210000000177000515000000000000000000;                                                                          // mov
      code[1233] = 'h00000023000000000000018c000015000000018b017516000000000001742100;                                                                          // moveLong
      code[1234] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1235] = 'h0000001f00000000000000000000010000000000006b20000000000000000000;                                                                          // label
      code[1236] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1237] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1238] = 'h000000220000000000000000018d210000000176000015000000000000000000;                                                                          // mov
      code[1239] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1240] = 'h0000002200000000000001770002150000000000017621000000000000000000;                                                                          // mov
      code[1241] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1242] = 'h0000002200000000000001670000150000000000017421000000000000000000;                                                                          // mov
      code[1243] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1244] = 'h000000220000000000000000018e210000000176000615000000000000000000;                                                                          // mov
      code[1245] = 'h000000220000000000000000018f21000000018e018d16000000000000000000;                                                                          // mov
      code[1246] = 'h0000001c000000000000001c0070210000000000018f21000000000001672100;                                                                          // jNe
      code[1247] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1248] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1249] = 'h0000002200000000000000000190210000000167000415000000000000000000;                                                                          // mov
      code[1250] = 'h0000002200000000000000000191210000000190017416000000000000000000;                                                                          // mov
      code[1251] = 'h0000002200000000000000000192210000000176000415000000000000000000;                                                                          // mov
      code[1252] = 'h000000220000000000000192018d160000000000019121000000000000000000;                                                                          // mov
      code[1253] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1254] = 'h0000002200000000000000000193210000000167000515000000000000000000;                                                                          // mov
      code[1255] = 'h0000002200000000000000000194210000000193017416000000000000000000;                                                                          // mov
      code[1256] = 'h0000002200000000000000000195210000000176000515000000000000000000;                                                                          // mov
      code[1257] = 'h000000220000000000000195018d160000000000019421000000000000000000;                                                                          // mov
      code[1258] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1259] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1260] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1261] = 'h0000002200000000000000000196210000000167000415000000000000000000;                                                                          // mov
      code[1262] = 'h0000003000000000000000000196210000000000017421000000000000062000;                                                                          // resize
      code[1263] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1264] = 'h0000000000000000000000000197210000000000018d21000000000000012000;                                                                          // add
      code[1265] = 'h0000002200000000000001760000150000000000019721000000000000000000;                                                                          // mov
      code[1266] = 'h0000002200000000000000000198210000000176000615000000000000000000;                                                                          // mov
      code[1267] = 'h0000002200000000000001980197160000000000017721000000000000000000;                                                                          // mov
      code[1268] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1269] = 'h0000002200000000000000000199210000000167000515000000000000000000;                                                                          // mov
      code[1270] = 'h0000003000000000000000000199210000000000017421000000000000072000;                                                                          // resize
      code[1271] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1272] = 'h0000001e00000000000000d00066210000000000000000000000000000000000;                                                                          // jmp
      code[1273] = 'h0000001e00000000000000260071210000000000000000000000000000000000;                                                                          // jmp
      code[1274] = 'h0000001f00000000000000000000010000000000007020000000000000000000;                                                                          // label
      code[1275] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1276] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1277] = 'h000000220000000000000000019a210000000167000415000000000000000000;                                                                          // mov
      code[1278] = 'h000000220000000000000000019b21000000019a017416000000000000000000;                                                                          // mov
      code[1279] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1280] = 'h000000220000000000000000019c210000000167000515000000000000000000;                                                                          // mov
      code[1281] = 'h000000220000000000000000019d21000000019c017416000000000000000000;                                                                          // mov
      code[1282] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1283] = 'h0000000e00000000000000000000010000000000017621000000000000002000;                                                                          // assertNe
      code[1284] = 'h000000220000000000000000019e210000000176000615000000000000000000;                                                                          // mov
      code[1285] = 'h000000050000000000000000019f210000000000019e21000000000001672100;                                                                          // arrayIndex
      code[1286] = 'h000000380000000000000000019f210000000000019f21000000000000012000;                                                                          // subtract
      code[1287] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1288] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1289] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1290] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1291] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1292] = 'h00000022000000000000000001a0210000000176000515000000000000000000;                                                                          // mov
      code[1293] = 'h0000003700000000000001a0019f160000000000019d21000000000000000000;                                                                          // shiftUp
      code[1294] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1295] = 'h00000022000000000000000001a1210000000176000615000000000000000000;                                                                          // mov
      code[1296] = 'h00000000000000000000000001a2210000000000019f21000000000000012000;                                                                          // add
      code[1297] = 'h0000003700000000000001a101a2160000000000017721000000000000000000;                                                                          // shiftUp
      code[1298] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1299] = 'h00000022000000000000000001a3210000000176000415000000000000000000;                                                                          // mov
      code[1300] = 'h0000003700000000000001a3019f160000000000019b21000000000000000000;                                                                          // shiftUp
      code[1301] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1302] = 'h0000000000000000000001760000150000000176000015000000000000012000;                                                                          // add
      code[1303] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1304] = 'h00000022000000000000000001a4210000000167000515000000000000000000;                                                                          // mov
      code[1305] = 'h00000030000000000000000001a4210000000000017421000000000000072000;                                                                          // resize
      code[1306] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1307] = 'h00000022000000000000000001a5210000000167000415000000000000000000;                                                                          // mov
      code[1308] = 'h00000030000000000000000001a5210000000000017421000000000000062000;                                                                          // resize
      code[1309] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1310] = 'h0000001e00000000000000aa0066210000000000000000000000000000000000;                                                                          // jmp
      code[1311] = 'h0000001f00000000000000000000010000000000007120000000000000000000;                                                                          // label
      code[1312] = 'h0000001f00000000000000000000010000000000006920000000000000000000;                                                                          // label
      code[1313] = 'h00000001000000000000000001a6210000000000000520000000000000000000;                                                                          // array
      code[1314] = 'h0000002200000000000001a60000150000000000017421000000000000000000;                                                                          // mov
      code[1315] = 'h0000002200000000000001a60002150000000000000020000000000000000000;                                                                          // mov
      code[1316] = 'h00000001000000000000000001a7210000000000000620000000000000000000;                                                                          // array
      code[1317] = 'h0000002200000000000001a6000415000000000001a721000000000000000000;                                                                          // mov
      code[1318] = 'h00000001000000000000000001a8210000000000000720000000000000000000;                                                                          // array
      code[1319] = 'h0000002200000000000001a6000515000000000001a821000000000000000000;                                                                          // mov
      code[1320] = 'h0000002200000000000001a60006150000000000000020000000000000000000;                                                                          // mov
      code[1321] = 'h0000002200000000000001a60003150000000000017221000000000000000000;                                                                          // mov
      code[1322] = 'h0000000000000000000001720001150000000172000115000000000000012000;                                                                          // add
      code[1323] = 'h0000002200000000000001a60001150000000172000115000000000000000000;                                                                          // mov
      code[1324] = 'h00000001000000000000000001a9210000000000000520000000000000000000;                                                                          // array
      code[1325] = 'h0000002200000000000001a90000150000000000017421000000000000000000;                                                                          // mov
      code[1326] = 'h0000002200000000000001a90002150000000000000020000000000000000000;                                                                          // mov
      code[1327] = 'h00000001000000000000000001aa210000000000000620000000000000000000;                                                                          // array
      code[1328] = 'h0000002200000000000001a9000415000000000001aa21000000000000000000;                                                                          // mov
      code[1329] = 'h00000001000000000000000001ab210000000000000720000000000000000000;                                                                          // array
      code[1330] = 'h0000002200000000000001a9000515000000000001ab21000000000000000000;                                                                          // mov
      code[1331] = 'h0000002200000000000001a90006150000000000000020000000000000000000;                                                                          // mov
      code[1332] = 'h0000002200000000000001a90003150000000000017221000000000000000000;                                                                          // mov
      code[1333] = 'h0000000000000000000001720001150000000172000115000000000000012000;                                                                          // add
      code[1334] = 'h0000002200000000000001a90001150000000172000115000000000000000000;                                                                          // mov
      code[1335] = 'h00000025000000000000000001ac210000000167000615000000000000000000;                                                                          // not
      code[1336] = 'h0000001c000000000000004c007221000000000001ac21000000000000002000;                                                                          // jNe
      code[1337] = 'h00000001000000000000000001ad210000000000000820000000000000000000;                                                                          // array
      code[1338] = 'h0000002200000000000001a6000615000000000001ad21000000000000000000;                                                                          // mov
      code[1339] = 'h00000001000000000000000001ae210000000000000820000000000000000000;                                                                          // array
      code[1340] = 'h0000002200000000000001a9000615000000000001ae21000000000000000000;                                                                          // mov
      code[1341] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1342] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1343] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1344] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1345] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1346] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1347] = 'h00000022000000000000000001af210000000167000415000000000000000000;                                                                          // mov
      code[1348] = 'h00000022000000000000000001b02100000001a9000415000000000000000000;                                                                          // mov
      code[1349] = 'h0000002300000000000001b000001500000001af017516000000000001742100;                                                                          // moveLong
      code[1350] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1351] = 'h00000022000000000000000001b1210000000167000515000000000000000000;                                                                          // mov
      code[1352] = 'h00000022000000000000000001b22100000001a9000515000000000000000000;                                                                          // mov
      code[1353] = 'h0000002300000000000001b200001500000001b1017516000000000001742100;                                                                          // moveLong
      code[1354] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1355] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1356] = 'h00000022000000000000000001b3210000000167000615000000000000000000;                                                                          // mov
      code[1357] = 'h00000022000000000000000001b42100000001a9000615000000000000000000;                                                                          // mov
      code[1358] = 'h00000000000000000000000001b5210000000000017421000000000000012000;                                                                          // add
      code[1359] = 'h0000002300000000000001b400001500000001b3017516000000000001b52100;                                                                          // moveLong
      code[1360] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1361] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1362] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1363] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1364] = 'h00000022000000000000000001b6210000000167000615000000000000000000;                                                                          // mov
      code[1365] = 'h00000022000000000000000001b72100000001a6000615000000000000000000;                                                                          // mov
      code[1366] = 'h00000000000000000000000001b8210000000000017421000000000000012000;                                                                          // add
      code[1367] = 'h0000002300000000000001b700001500000001b6000015000000000001b82100;                                                                          // moveLong
      code[1368] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1369] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1370] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1371] = 'h00000022000000000000000001b9210000000167000415000000000000000000;                                                                          // mov
      code[1372] = 'h00000022000000000000000001ba2100000001a6000415000000000000000000;                                                                          // mov
      code[1373] = 'h0000002300000000000001ba00001500000001b9000015000000000001742100;                                                                          // moveLong
      code[1374] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1375] = 'h00000022000000000000000001bb210000000167000515000000000000000000;                                                                          // mov
      code[1376] = 'h00000022000000000000000001bc2100000001a6000515000000000000000000;                                                                          // mov
      code[1377] = 'h0000002300000000000001bc00001500000001bb000015000000000001742100;                                                                          // moveLong
      code[1378] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1379] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1380] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1381] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1382] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1383] = 'h00000022000000000000000001bd2100000001a6000015000000000000000000;                                                                          // mov
      code[1384] = 'h00000000000000000000000001be21000000000001bd21000000000000012000;                                                                          // add
      code[1385] = 'h00000022000000000000000001bf2100000001a6000615000000000000000000;                                                                          // mov
      code[1386] = 'h0000001f00000000000000000000010000000000007420000000000000000000;                                                                          // label
      code[1387] = 'h00000022000000000000000001c0210000000000000020000000000000000000;                                                                          // mov
      code[1388] = 'h0000001f00000000000000000000010000000000007520000000000000000000;                                                                          // label
      code[1389] = 'h000000180000000000000006007721000000000001c021000000000001be2100;                                                                          // jGe
      code[1390] = 'h00000022000000000000000001c12100000001bf01c016000000000000000000;                                                                          // mov
      code[1391] = 'h0000002200000000000001c1000215000000000001a621000000000000000000;                                                                          // mov
      code[1392] = 'h0000001f00000000000000000000010000000000007620000000000000000000;                                                                          // label
      code[1393] = 'h00000000000000000000000001c021000000000001c021000000000000012000;                                                                          // add
      code[1394] = 'h0000001e00000000fffffffa0075210000000000000000000000000000000000;                                                                          // jmp
      code[1395] = 'h0000001f00000000000000000000010000000000007720000000000000000000;                                                                          // label
      code[1396] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1397] = 'h00000022000000000000000001c22100000001a9000015000000000000000000;                                                                          // mov
      code[1398] = 'h00000000000000000000000001c321000000000001c221000000000000012000;                                                                          // add
      code[1399] = 'h00000022000000000000000001c42100000001a9000615000000000000000000;                                                                          // mov
      code[1400] = 'h0000001f00000000000000000000010000000000007820000000000000000000;                                                                          // label
      code[1401] = 'h00000022000000000000000001c5210000000000000020000000000000000000;                                                                          // mov
      code[1402] = 'h0000001f00000000000000000000010000000000007920000000000000000000;                                                                          // label
      code[1403] = 'h000000180000000000000006007b21000000000001c521000000000001c32100;                                                                          // jGe
      code[1404] = 'h00000022000000000000000001c62100000001c401c516000000000000000000;                                                                          // mov
      code[1405] = 'h0000002200000000000001c6000215000000000001a921000000000000000000;                                                                          // mov
      code[1406] = 'h0000001f00000000000000000000010000000000007a20000000000000000000;                                                                          // label
      code[1407] = 'h00000000000000000000000001c521000000000001c521000000000000012000;                                                                          // add
      code[1408] = 'h0000001e00000000fffffffa0079210000000000000000000000000000000000;                                                                          // jmp
      code[1409] = 'h0000001f00000000000000000000010000000000007b20000000000000000000;                                                                          // label
      code[1410] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1411] = 'h0000001e000000000000001d0073210000000000000000000000000000000000;                                                                          // jmp
      code[1412] = 'h0000001f00000000000000000000010000000000007220000000000000000000;                                                                          // label
      code[1413] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1414] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1415] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1416] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1417] = 'h00000022000000000000000001c7210000000167000515000000000000000000;                                                                          // mov
      code[1418] = 'h00000022000000000000000001c82100000001a6000515000000000000000000;                                                                          // mov
      code[1419] = 'h0000002300000000000001c800001500000001c7000015000000000001742100;                                                                          // moveLong
      code[1420] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1421] = 'h00000022000000000000000001c9210000000167000415000000000000000000;                                                                          // mov
      code[1422] = 'h00000022000000000000000001ca2100000001a6000415000000000000000000;                                                                          // mov
      code[1423] = 'h0000002300000000000001ca00001500000001c9000015000000000001742100;                                                                          // moveLong
      code[1424] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1425] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1426] = 'h00000001000000000000000001cb210000000000000820000000000000000000;                                                                          // array
      code[1427] = 'h000000220000000000000167000615000000000001cb21000000000000000000;                                                                          // mov
      code[1428] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1429] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1430] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1431] = 'h00000022000000000000000001cc210000000167000415000000000000000000;                                                                          // mov
      code[1432] = 'h00000022000000000000000001cd2100000001a9000415000000000000000000;                                                                          // mov
      code[1433] = 'h0000002300000000000001cd00001500000001cc017516000000000001742100;                                                                          // moveLong
      code[1434] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1435] = 'h00000022000000000000000001ce210000000167000515000000000000000000;                                                                          // mov
      code[1436] = 'h00000022000000000000000001cf2100000001a9000515000000000000000000;                                                                          // mov
      code[1437] = 'h0000002300000000000001cf00001500000001ce017516000000000001742100;                                                                          // moveLong
      code[1438] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1439] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1440] = 'h0000001f00000000000000000000010000000000007320000000000000000000;                                                                          // label
      code[1441] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1442] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1443] = 'h00000022000000000000000001d0210000000167000515000000000000000000;                                                                          // mov
      code[1444] = 'h00000022000000000000000001d12100000001d0017416000000000000000000;                                                                          // mov
      code[1445] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1446] = 'h0000002200000000000001a90002150000000000016721000000000000000000;                                                                          // mov
      code[1447] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1448] = 'h00000022000000000000000001d2210000000167000415000000000000000000;                                                                          // mov
      code[1449] = 'h00000022000000000000000001d32100000001d2017416000000000000000000;                                                                          // mov
      code[1450] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1451] = 'h0000002200000000000001a60002150000000000016721000000000000000000;                                                                          // mov
      code[1452] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1453] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1454] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1455] = 'h00000022000000000000000001d4210000000167000515000000000000000000;                                                                          // mov
      code[1456] = 'h00000030000000000000000001d4210000000000000120000000000000072000;                                                                          // resize
      code[1457] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1458] = 'h00000022000000000000000001d5210000000167000615000000000000000000;                                                                          // mov
      code[1459] = 'h0000002200000000000001d5000015000000000001a621000000000000000000;                                                                          // mov
      code[1460] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1461] = 'h0000002200000000000001670000150000000000000120000000000000000000;                                                                          // mov
      code[1462] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1463] = 'h00000022000000000000000001d6210000000167000415000000000000000000;                                                                          // mov
      code[1464] = 'h00000030000000000000000001d6210000000000000120000000000000062000;                                                                          // resize
      code[1465] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1466] = 'h00000022000000000000000001d7210000000167000515000000000000000000;                                                                          // mov
      code[1467] = 'h0000002200000000000001d7000015000000000001d121000000000000000000;                                                                          // mov
      code[1468] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1469] = 'h00000022000000000000000001d8210000000167000615000000000000000000;                                                                          // mov
      code[1470] = 'h00000030000000000000000001d8210000000000000220000000000000082000;                                                                          // resize
      code[1471] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1472] = 'h00000022000000000000000001d9210000000167000415000000000000000000;                                                                          // mov
      code[1473] = 'h0000002200000000000001d9000015000000000001d321000000000000000000;                                                                          // mov
      code[1474] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1475] = 'h00000022000000000000000001da210000000167000615000000000000000000;                                                                          // mov
      code[1476] = 'h0000002200000000000001da000115000000000001a921000000000000000000;                                                                          // mov
      code[1477] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1478] = 'h0000001e00000000000000020066210000000000000000000000000000000000;                                                                          // jmp
      code[1479] = 'h0000001e00000000000000060068210000000000000000000000000000000000;                                                                          // jmp
      code[1480] = 'h0000001f00000000000000000000010000000000006620000000000000000000;                                                                          // label
      code[1481] = 'h0000002200000000000000000170210000000000000120000000000000000000;                                                                          // mov
      code[1482] = 'h0000001e00000000000000030068210000000000000000000000000000000000;                                                                          // jmp
      code[1483] = 'h0000001f00000000000000000000010000000000006720000000000000000000;                                                                          // label
      code[1484] = 'h0000002200000000000000000170210000000000000020000000000000000000;                                                                          // mov
      code[1485] = 'h0000001f00000000000000000000010000000000006820000000000000000000;                                                                          // label
      code[1486] = 'h0000001f00000000000000000000010000000000000620000000000000000000;                                                                          // label
      code[1487] = 'h0000001f00000000000000000000010000000000000720000000000000000000;                                                                          // label
      code[1488] = 'h0000001f00000000000000000000010000000000000820000000000000000000;                                                                          // label
      code[1489] = 'h0000001300000000000000000003210000000000000420000000000000000000;                                                                          // free
      code[1490] = 'h0000001f00000000000000000000010000000000000320000000000000000000;                                                                          // label
      code[1491] = 'h0000003800000000000000000001210000000000000121000000000000012000;                                                                          // subtract
      code[1492] = 'h0000001e00000000fffffa3a0002210000000000000000000000000000000000;                                                                          // jmp
      code[1493] = 'h0000001f00000000000000000000010000000000000420000000000000000000;                                                                          // label
      code[1494] = 'h00000022000000000000000001db210000000000000120000000000000000000;                                                                          // mov
      code[1495] = 'h00000035000000000000000001db210000000000001f20000000000000000000;                                                                          // shiftLeft
      code[1496] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1497] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1498] = 'h00000001000000000000000001dc210000000000000420000000000000000000;                                                                          // array
      code[1499] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1500] = 'h00000022000000000000000001dd210000000000000315000000000000000000;                                                                          // mov
      code[1501] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1502] = 'h00000001000000000000000001de210000000000000420000000000000000000;                                                                          // array
      code[1503] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1504] = 'h0000001c0000000000000009007c21000000000001dd21000000000000002000;                                                                          // jNe
      code[1505] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1506] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1507] = 'h0000002200000000000001de0001150000000000000320000000000000000000;                                                                          // mov
      code[1508] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1509] = 'h0000002200000000000001de000015000000000001dd21000000000000000000;                                                                          // mov
      code[1510] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1511] = 'h0000002200000000000001de0002150000000000000020000000000000000000;                                                                          // mov
      code[1512] = 'h0000001e0000000000000016007d210000000000000000000000000000000000;                                                                          // jmp
      code[1513] = 'h0000001f00000000000000000000010000000000007c20000000000000000000;                                                                          // label
      code[1514] = 'h0000001f00000000000000000000010000000000007e20000000000000000000;                                                                          // label
      code[1515] = 'h00000022000000000000000001df210000000000000020000000000000000000;                                                                          // mov
      code[1516] = 'h0000001f00000000000000000000010000000000007f20000000000000000000;                                                                          // label
      code[1517] = 'h000000180000000000000009008121000000000001df21000000000000632000;                                                                          // jGe
      code[1518] = 'h00000025000000000000000001e02100000001dd000615000000000000000000;                                                                          // not
      code[1519] = 'h0000001d0000000000000007008121000000000001e021000000000000000000;                                                                          // jTrue
      code[1520] = 'h00000022000000000000000001e12100000001dd000615000000000000000000;                                                                          // mov
      code[1521] = 'h00000022000000000000000001e22100000001e1000015000000000000000000;                                                                          // mov
      code[1522] = 'h00000022000000000000000001dd21000000000001e221000000000000000000;                                                                          // mov
      code[1523] = 'h0000001f00000000000000000000010000000000008020000000000000000000;                                                                          // label
      code[1524] = 'h00000000000000000000000001df21000000000001df21000000000000012000;                                                                          // add
      code[1525] = 'h0000001e00000000fffffff7007f210000000000000000000000000000000000;                                                                          // jmp
      code[1526] = 'h0000001f00000000000000000000010000000000008120000000000000000000;                                                                          // label
      code[1527] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1528] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1529] = 'h0000002200000000000001de0001150000000000000120000000000000000000;                                                                          // mov
      code[1530] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1531] = 'h0000002200000000000001de000015000000000001dd21000000000000000000;                                                                          // mov
      code[1532] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1533] = 'h0000002200000000000001de0002150000000000000020000000000000000000;                                                                          // mov
      code[1534] = 'h0000001f00000000000000000000010000000000007d20000000000000000000;                                                                          // label
      code[1535] = 'h0000001f00000000000000000000010000000000008220000000000000000000;                                                                          // label
      code[1536] = 'h00000022000000000000000001e32100000001de000115000000000000000000;                                                                          // mov
      code[1537] = 'h00000016000000000000006f008521000000000001e321000000000000032000;                                                                          // jEq
      code[1538] = 'h0000002300000000000001dc00001500000001de000015000000000000032000;                                                                          // moveLong
      code[1539] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1540] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1541] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1542] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1543] = 'h00000022000000000000000001e42100000001dc000015000000000000000000;                                                                          // mov
      code[1544] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1545] = 'h00000022000000000000000001e52100000001dc000215000000000000000000;                                                                          // mov
      code[1546] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1547] = 'h00000022000000000000000001e62100000001e4000415000000000000000000;                                                                          // mov
      code[1548] = 'h00000022000000000000000001e72100000001e601e516000000000000000000;                                                                          // mov
      code[1549] = 'h000000260000000000000000000001000000000001e721000000000000000000;                                                                          // out
      code[1550] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1551] = 'h0000001f00000000000000000000010000000000008620000000000000000000;                                                                          // label
      code[1552] = 'h00000022000000000000000001e82100000001de000015000000000000000000;                                                                          // mov
      code[1553] = 'h00000025000000000000000001e92100000001e8000615000000000000000000;                                                                          // not
      code[1554] = 'h000000160000000000000034008a21000000000001e921000000000000002000;                                                                          // jEq
      code[1555] = 'h00000000000000000000000001ea2100000001de000215000000000000012000;                                                                          // add
      code[1556] = 'h00000022000000000000000001eb2100000001e8000015000000000000000000;                                                                          // mov
      code[1557] = 'h000000180000000000000009008b21000000000001ea21000000000001eb2100;                                                                          // jGe
      code[1558] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1559] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1560] = 'h0000002200000000000001de0001150000000000000120000000000000000000;                                                                          // mov
      code[1561] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1562] = 'h0000002200000000000001de000015000000000001e821000000000000000000;                                                                          // mov
      code[1563] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1564] = 'h0000002200000000000001de000215000000000001ea21000000000000000000;                                                                          // mov
      code[1565] = 'h0000001e000000000000004e0089210000000000000000000000000000000000;                                                                          // jmp
      code[1566] = 'h0000001f00000000000000000000010000000000008b20000000000000000000;                                                                          // label
      code[1567] = 'h00000022000000000000000001ec2100000001e8000215000000000000000000;                                                                          // mov
      code[1568] = 'h00000016000000000000001d008c21000000000001ec21000000000000002000;                                                                          // jEq
      code[1569] = 'h0000001f00000000000000000000010000000000008d20000000000000000000;                                                                          // label
      code[1570] = 'h00000022000000000000000001ed210000000000000020000000000000000000;                                                                          // mov
      code[1571] = 'h0000001f00000000000000000000010000000000008e20000000000000000000;                                                                          // label
      code[1572] = 'h000000180000000000000018009021000000000001ed21000000000000632000;                                                                          // jGe
      code[1573] = 'h00000022000000000000000001ee2100000001ec000015000000000000000000;                                                                          // mov
      code[1574] = 'h0000000e0000000000000000000001000000000001ec21000000000000002000;                                                                          // assertNe
      code[1575] = 'h00000022000000000000000001ef2100000001ec000615000000000000000000;                                                                          // mov
      code[1576] = 'h00000005000000000000000001f021000000000001ef21000000000001e82100;                                                                          // arrayIndex
      code[1577] = 'h00000038000000000000000001f021000000000001f021000000000000012000;                                                                          // subtract
      code[1578] = 'h0000001c0000000000000005009121000000000001f021000000000001ee2100;                                                                          // jNe
      code[1579] = 'h00000022000000000000000001e821000000000001ec21000000000000000000;                                                                          // mov
      code[1580] = 'h00000022000000000000000001ec2100000001e8000215000000000000000000;                                                                          // mov
      code[1581] = 'h00000017000000000000000f009021000000000001ec21000000000000000000;                                                                          // jFalse
      code[1582] = 'h0000001e000000000000000a0092210000000000000000000000000000000000;                                                                          // jmp
      code[1583] = 'h0000001f00000000000000000000010000000000009120000000000000000000;                                                                          // label
      code[1584] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1585] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1586] = 'h0000002200000000000001de000015000000000001ec21000000000000000000;                                                                          // mov
      code[1587] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1588] = 'h0000002200000000000001de0001150000000000000120000000000000000000;                                                                          // mov
      code[1589] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1590] = 'h0000002200000000000001de000215000000000001f021000000000000000000;                                                                          // mov
      code[1591] = 'h0000001e00000000000000340089210000000000000000000000000000000000;                                                                          // jmp
      code[1592] = 'h0000001f00000000000000000000010000000000009220000000000000000000;                                                                          // label
      code[1593] = 'h0000001f00000000000000000000010000000000008f20000000000000000000;                                                                          // label
      code[1594] = 'h00000000000000000000000001ed21000000000001ed21000000000000012000;                                                                          // add
      code[1595] = 'h0000001e00000000ffffffe8008e210000000000000000000000000000000000;                                                                          // jmp
      code[1596] = 'h0000001f00000000000000000000010000000000009020000000000000000000;                                                                          // label
      code[1597] = 'h0000001f00000000000000000000010000000000008c20000000000000000000;                                                                          // label
      code[1598] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1599] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1600] = 'h0000002200000000000001de0001150000000000000320000000000000000000;                                                                          // mov
      code[1601] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1602] = 'h0000002200000000000001de000015000000000001e821000000000000000000;                                                                          // mov
      code[1603] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1604] = 'h0000002200000000000001de0002150000000000000020000000000000000000;                                                                          // mov
      code[1605] = 'h0000001e00000000000000260089210000000000000000000000000000000000;                                                                          // jmp
      code[1606] = 'h0000001f00000000000000000000010000000000008a20000000000000000000;                                                                          // label
      code[1607] = 'h00000000000000000000000001f12100000001de000215000000000000012000;                                                                          // add
      code[1608] = 'h00000022000000000000000001f22100000001e8000615000000000000000000;                                                                          // mov
      code[1609] = 'h00000022000000000000000001f32100000001f201f116000000000000000000;                                                                          // mov
      code[1610] = 'h0000001c0000000000000009009321000000000001f321000000000000002000;                                                                          // jNe
      code[1611] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1612] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1613] = 'h0000002200000000000001de000015000000000001f321000000000000000000;                                                                          // mov
      code[1614] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1615] = 'h0000002200000000000001de0001150000000000000320000000000000000000;                                                                          // mov
      code[1616] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1617] = 'h0000002200000000000001de0002150000000000000020000000000000000000;                                                                          // mov
      code[1618] = 'h0000001e00000000000000160094210000000000000000000000000000000000;                                                                          // jmp
      code[1619] = 'h0000001f00000000000000000000010000000000009320000000000000000000;                                                                          // label
      code[1620] = 'h0000001f00000000000000000000010000000000009520000000000000000000;                                                                          // label
      code[1621] = 'h00000022000000000000000001f4210000000000000020000000000000000000;                                                                          // mov
      code[1622] = 'h0000001f00000000000000000000010000000000009620000000000000000000;                                                                          // label
      code[1623] = 'h000000180000000000000009009821000000000001f421000000000000632000;                                                                          // jGe
      code[1624] = 'h00000025000000000000000001f52100000001f3000615000000000000000000;                                                                          // not
      code[1625] = 'h0000001d0000000000000007009821000000000001f521000000000000000000;                                                                          // jTrue
      code[1626] = 'h00000022000000000000000001f62100000001f3000615000000000000000000;                                                                          // mov
      code[1627] = 'h00000022000000000000000001f72100000001f6000015000000000000000000;                                                                          // mov
      code[1628] = 'h00000022000000000000000001f321000000000001f721000000000000000000;                                                                          // mov
      code[1629] = 'h0000001f00000000000000000000010000000000009720000000000000000000;                                                                          // label
      code[1630] = 'h00000000000000000000000001f421000000000001f421000000000000012000;                                                                          // add
      code[1631] = 'h0000001e00000000fffffff70096210000000000000000000000000000000000;                                                                          // jmp
      code[1632] = 'h0000001f00000000000000000000010000000000009820000000000000000000;                                                                          // label
      code[1633] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1634] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1635] = 'h0000002200000000000001de000015000000000001f321000000000000000000;                                                                          // mov
      code[1636] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1637] = 'h0000002200000000000001de0001150000000000000120000000000000000000;                                                                          // mov
      code[1638] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1639] = 'h0000002200000000000001de0002150000000000000020000000000000000000;                                                                          // mov
      code[1640] = 'h0000001f00000000000000000000010000000000009420000000000000000000;                                                                          // label
      code[1641] = 'h0000001f00000000000000000000010000000000008720000000000000000000;                                                                          // label
      code[1642] = 'h0000001f00000000000000000000010000000000008820000000000000000000;                                                                          // label
      code[1643] = 'h0000001f00000000000000000000010000000000008920000000000000000000;                                                                          // label
      code[1644] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
      code[1645] = 'h0000001e00000000ffffff920082210000000000000000000000000000000000;                                                                          // jmp
      code[1646] = 'h0000001f00000000000000000000010000000000008320000000000000000000;                                                                          // label
      code[1647] = 'h0000001f00000000000000000000010000000000008420000000000000000000;                                                                          // label
      code[1648] = 'h0000001f00000000000000000000010000000000008520000000000000000000;                                                                          // label
      code[1649] = 'h0000002800000000000000000000010000000000000000000000000000000000;                                                                          // parallelStart
      code[1650] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1651] = 'h00000013000000000000000001dc210000000000000420000000000000000000;                                                                          // free
      code[1652] = 'h0000002700000000000000000000010000000000000000000000000000000000;                                                                          // parallelContinue
      code[1653] = 'h00000013000000000000000001de210000000000000420000000000000000000;                                                                          // free
      code[1654] = 'h0000002900000000000000000000010000000000000000000000000000000000;                                                                          // parallelStop
    end
  endtask
                                                                                // Load program 'In_test' into code memory
  task In_test();
    begin
      NInstructionEnd = 9;
      code[   0] = 'h0000001f00000000000000000000010000000000000120000000000000000000;                                                                          // label
      code[   1] = 'h0000001500000000000000000000210000000000000000000000000000000000;                                                                          // inSize
      code[   2] = 'h0000001700000000000000060003210000000000000021000000000000000000;                                                                          // jFalse
      code[   3] = 'h0000001400000000000000000001210000000000000000000000000000000000;                                                                          // in
      code[   4] = 'h0000002600000000000000000000010000000000000021000000000000000000;                                                                          // out
      code[   5] = 'h0000002600000000000000000000010000000000000121000000000000000000;                                                                          // out
      code[   6] = 'h0000001f00000000000000000000010000000000000220000000000000000000;                                                                          // label
      code[   7] = 'h0000001e00000000fffffff90001210000000000000000000000000000000000;                                                                          // jmp
      code[   8] = 'h0000001f00000000000000000000010000000000000320000000000000000000;                                                                          // label
    end
  endtask

//Memory access functions for instruction execution

  task setMemory();                                                             // Set the target memory location updating the containing array size if necessary
    begin
      case(targetArena)
        1: fork                                                                 // Update array
          heapMem[targetLocation] = result;
          arraySizes[targetLocationArea]  =
          arraySizes[targetLocationArea] >  targetIndex ?
          arraySizes[targetLocationArea]  : targetIndex + 1;
        join
        2: localMem[targetLocation] = result;                                   // Local memory
      endcase
    end
  endtask

//Implementation of each instruction

  task add_instruction();                                                       // Add
    begin
      result = source1Value + source2Value;
      setMemory();
    end
  endtask

  task array_instruction();                                                     // Array
    begin
      if (freedArraysTop > 0) begin                                             // Reuse an array
        result = freedArrays[--freedArraysTop];
      end
      else begin
        result = allocs++;                                                      // Array zero means undefined
      end

      arraySizes[targetLocationArea] = 0;                                       // Zero array length
      setMemory();                                                              // Save address of array
    end
  endtask

  task free_instruction();
    begin                                                                       // Free
      freedArrays[freedArraysTop++] = targetValue;
      arraySizes[targetValue] = 0;                                              // Zero array length
    end
  endtask

  task mov_instruction();                                                       // Mov
    begin
      result = source1Value;
      //$display("%4d = Mov %d(%d), %d", result, targetLocation, targetArena, source1Value);
      setMemory();                                                              // Save result in target
    end
  endtask


  task not_instruction();                                                       // Not
    begin
      result = source1Value ? 0 : 1;
      setMemory();                                                              // Save result in target
    end
  endtask

  task resize_instruction();                                                    // Resize
    begin
      result = source1Value;
      p = localMem[targetLocation];
      fork
        heapMem[p * NArea] = result;
        q = heapMem[p * NArea];
      join
    end
  endtask

  task subtract_instruction();                                                  // Subtract
    begin
      result = source1Value - source2Value;
      setMemory();                                                              // Save result in target
    end
  endtask

  task out_instruction();                                                       // Out
    begin
//$display("AAAAA %d",source1Value);
      outMem[outMemPos++] = source1Value;
    end
  endtask

  task arrayIndex_instruction();
    begin                                                                       // ArrayIndex
      fork
        q = source1Value * NArea;                                               // Array location
        p = arraySizes[source1Value];                                           // Length of array
        result = 0;
      join
      case(p)                                                                   // Arrays can be dynamic but only up to a fixed size so that we can unroll the loop that finds an element
        1:
            begin if (heapMem[q+0] == source2Value) result = 1; end
        2:
          fork
            begin if (heapMem[q+0] == source2Value) result = 1; end
            begin if (heapMem[q+1] == source2Value) result = 2; end
          join
        3:
          fork
            begin if (heapMem[q+0] == source2Value) result = 1; end
            begin if (heapMem[q+1] == source2Value) result = 2; end
            begin if (heapMem[q+2] == source2Value) result = 3; end
          join
        4:
          fork
            begin if (heapMem[q+0] == source2Value) result = 1; end
            begin if (heapMem[q+1] == source2Value) result = 2; end
            begin if (heapMem[q+2] == source2Value) result = 3; end
            begin if (heapMem[q+3] == source2Value) result = 4; end
          join
        5:
          fork
            begin if (heapMem[q+0] == source2Value) result = 1; end
            begin if (heapMem[q+1] == source2Value) result = 2; end
            begin if (heapMem[q+2] == source2Value) result = 3; end
            begin if (heapMem[q+3] == source2Value) result = 4; end
            begin if (heapMem[q+4] == source2Value) result = 5; end
          join
        6:
          fork
            begin if (heapMem[q+0] == source2Value) result = 1; end
            begin if (heapMem[q+1] == source2Value) result = 2; end
            begin if (heapMem[q+2] == source2Value) result = 3; end
            begin if (heapMem[q+3] == source2Value) result = 4; end
            begin if (heapMem[q+4] == source2Value) result = 5; end
            begin if (heapMem[q+5] == source2Value) result = 6; end
          join
        7:
          fork
            begin if (heapMem[q+0] == source2Value) result = 1; end
            begin if (heapMem[q+1] == source2Value) result = 2; end
            begin if (heapMem[q+2] == source2Value) result = 3; end
            begin if (heapMem[q+3] == source2Value) result = 4; end
            begin if (heapMem[q+4] == source2Value) result = 5; end
            begin if (heapMem[q+5] == source2Value) result = 6; end
            begin if (heapMem[q+6] == source2Value) result = 7; end
          join
      endcase
      setMemory();
    end
  endtask

  task arrayCountGreater_instruction();
    begin                                                                       // ArrayIndex
      fork
        q = source1Value * NArea;                                               // Array location
        p = arraySizes[source1Value];                                           // Length of array
        result = 0;
        r1 = 0; r2 = 0; r3 = 0; r4 = 0; r5 = 0; r6 = 0; r7 = 0; r8 = 0;
      join;
      case(p)                                                                   // Arrays can be dynamic but only up to a fixed size so that we can unroll the loop that finds an element
        1:
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
        2:
          fork
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
            begin if (heapMem[q+1] > source2Value) r2 = 1; end
          join
        3:
          fork
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
            begin if (heapMem[q+1] > source2Value) r2 = 1; end
            begin if (heapMem[q+2] > source2Value) r3 = 1; end
          join
        4:
          fork
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
            begin if (heapMem[q+1] > source2Value) r2 = 1; end
            begin if (heapMem[q+2] > source2Value) r3 = 1; end
            begin if (heapMem[q+3] > source2Value) r4 = 1; end
          join
        5:
          fork
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
            begin if (heapMem[q+1] > source2Value) r2 = 1; end
            begin if (heapMem[q+2] > source2Value) r3 = 1; end
            begin if (heapMem[q+3] > source2Value) r4 = 1; end
            begin if (heapMem[q+4] > source2Value) r5 = 1; end
          join
        6:
          fork
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
            begin if (heapMem[q+1] > source2Value) r2 = 1; end
            begin if (heapMem[q+2] > source2Value) r3 = 1; end
            begin if (heapMem[q+3] > source2Value) r4 = 1; end
            begin if (heapMem[q+4] > source2Value) r5 = 1; end
            begin if (heapMem[q+5] > source2Value) r6 = 1; end
          join
        7:
          fork
            begin if (heapMem[q+0] > source2Value) r1 = 1; end
            begin if (heapMem[q+1] > source2Value) r2 = 1; end
            begin if (heapMem[q+2] > source2Value) r3 = 1; end
            begin if (heapMem[q+3] > source2Value) r4 = 1; end
            begin if (heapMem[q+4] > source2Value) r5 = 1; end
            begin if (heapMem[q+5] > source2Value) r6 = 1; end
            begin if (heapMem[q+6] > source2Value) r7 = 1; end
          join
      endcase
      result = r1 + r2 + r3 + r4 + r5 + r6 + r7 + r8;
      setMemory();
    end
  endtask

  task arrayCountLess_instruction();
    begin                                                                       // ArrayIndex
      fork
        q = source1Value * NArea;                                               // Array location
        p = arraySizes[source1Value];                                           // Length of array
        result = 0;
        r1 = 0; r2 = 0; r3 = 0; r4 = 0; r5 = 0; r6 = 0; r7 = 0; r8 = 0;
      join
      case(p)                                                                   // Arrays can be dynamic but only up to a fixed size so that we can unroll the loop that finds an element
        1:
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
        2:
          fork
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
            begin if (heapMem[q+1] < source2Value) r2 = 1; end
          join
        3:
          fork
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
            begin if (heapMem[q+1] < source2Value) r2 = 1; end
            begin if (heapMem[q+2] < source2Value) r3 = 1; end
          join
        4:
          fork
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
            begin if (heapMem[q+1] < source2Value) r2 = 1; end
            begin if (heapMem[q+2] < source2Value) r3 = 1; end
            begin if (heapMem[q+3] < source2Value) r4 = 1; end
          join
        5:
          fork
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
            begin if (heapMem[q+1] < source2Value) r2 = 1; end
            begin if (heapMem[q+2] < source2Value) r3 = 1; end
            begin if (heapMem[q+3] < source2Value) r4 = 1; end
            begin if (heapMem[q+4] < source2Value) r5 = 1; end
          join
        6:
          fork
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
            begin if (heapMem[q+1] < source2Value) r2 = 1; end
            begin if (heapMem[q+2] < source2Value) r3 = 1; end
            begin if (heapMem[q+3] < source2Value) r4 = 1; end
            begin if (heapMem[q+4] < source2Value) r5 = 1; end
            begin if (heapMem[q+5] < source2Value) r6 = 1; end
          join
        7:
          fork
            begin if (heapMem[q+0] < source2Value) r1 = 1; end
            begin if (heapMem[q+1] < source2Value) r2 = 1; end
            begin if (heapMem[q+2] < source2Value) r3 = 1; end
            begin if (heapMem[q+3] < source2Value) r4 = 1; end
            begin if (heapMem[q+4] < source2Value) r5 = 1; end
            begin if (heapMem[q+5] < source2Value) r6 = 1; end
            begin if (heapMem[q+6] < source2Value) r7 = 1; end
          join
      endcase
      result = r1 + r2 + r3 + r4 + r5 + r6 + r7 + r8;
      setMemory();
    end
  endtask

  task shiftLeft_instruction();
    begin                                                                       // shiftLeft
      result = targetValue << source1Value;
      setMemory();
    end
  endtask

  task shiftRight_instruction();
    begin                                                                       // shiftLeft
      result = targetValue >> source1Value;
      setMemory();
    end
  endtask

  task jEq_instruction();
    begin                                                                       // Jeq
      if (source1Value == source2Value) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jFalse_instruction();
    begin                                                                       // jFalse
      if (source1Value == 0) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jGe_instruction();
    begin                                                                       // jGe
      if (source1Value >= source2Value) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jGt_instruction();
    begin                                                                       // jGt
      if (source1Value >  source2Value) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jLe_instruction();
    begin                                                                       // jLe
      if (source1Value <= source2Value) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jLt_instruction();
    begin                                                                       // jLt
      if (source1Value <  source2Value) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jNe_instruction();
    begin                                                                       // jNe
      if (source1Value != source2Value) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jTrue_instruction();
    begin                                                                       // jTrue
      if (source1Value != 0) begin
        ip += targetArea - 1;
      end
    end
  endtask

  task jmp_instruction();
    begin                                                                       // jmp
      ip += targetArea - 1;
    end
  endtask

  task push_instruction();                                                      // push
    begin
      p = arraySizes[targetValue];
      if (p + 1 < NArea) begin
        heapMem[p] = source1Value;
        arraySizes[targetValue] = p + 1;
        result = source1Value;
      end
    end
  endtask

  task pop_instruction();                                                       // pop
    begin
      p = arraySizes[source1Value];
      if (p > 0) begin
        p--;
        arraySizes[source1Value] = p;
        result = heapMem[p];
        setMemory();
        result = source1Value;
      end
    end
  endtask

  task arraySize_instruction();
    begin                                                                       // arraySize
      result = arraySizes[source1Value];
      setMemory();
    end
  endtask
                                                                                // Shift up an array in parallel by first copying every element in parallel then copying back just the elements we need into their new positions
  task shiftUp_instruction();
    begin
      if (targetIndex < NArea) begin
        p = targetLocationArea * NArea;                                         // Array Start
        fork
          arraySizes[targetLocationArea] = arraySizes[targetLocationArea] + 1;  // New size of array
          if (NArea > 0) arrayShift[0] = heapMem[p + 0];                        // Move data into staging area
          if (NArea > 1) arrayShift[1] = heapMem[p + 1];
          if (NArea > 2) arrayShift[2] = heapMem[p + 2];
          if (NArea > 3) arrayShift[3] = heapMem[p + 3];
          if (NArea > 4) arrayShift[4] = heapMem[p + 4];
          if (NArea > 5) arrayShift[5] = heapMem[p + 5];
          if (NArea > 6) arrayShift[6] = heapMem[p + 6];
          if (NArea > 7) arrayShift[7] = heapMem[p + 7];
          if (NArea > 8) arrayShift[8] = heapMem[p + 8];
          if (NArea > 9) arrayShift[9] = heapMem[p + 9];
        join
        case(targetIndex)                                                       // Destage data into one position higher
          0: fork
            if (NArea > 0) heapMem[p + 0] = source1Value;
            if (NArea > 1) heapMem[p + 1] = arrayShift[0];
            if (NArea > 2) heapMem[p + 2] = arrayShift[1];
            if (NArea > 3) heapMem[p + 3] = arrayShift[2];
            if (NArea > 4) heapMem[p + 4] = arrayShift[3];
            if (NArea > 5) heapMem[p + 5] = arrayShift[4];
            if (NArea > 6) heapMem[p + 6] = arrayShift[5];
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          1: fork
            if (NArea > 1) heapMem[p + 1] = source1Value;
            if (NArea > 2) heapMem[p + 2] = arrayShift[1];
            if (NArea > 3) heapMem[p + 3] = arrayShift[2];
            if (NArea > 4) heapMem[p + 4] = arrayShift[3];
            if (NArea > 5) heapMem[p + 5] = arrayShift[4];
            if (NArea > 6) heapMem[p + 6] = arrayShift[5];
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          2: fork
            if (NArea > 2) heapMem[p + 2] = source1Value;
            if (NArea > 3) heapMem[p + 3] = arrayShift[2];
            if (NArea > 4) heapMem[p + 4] = arrayShift[3];
            if (NArea > 5) heapMem[p + 5] = arrayShift[4];
            if (NArea > 6) heapMem[p + 6] = arrayShift[5];
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          3: fork
            if (NArea > 3) heapMem[p + 3] = source1Value;
            if (NArea > 4) heapMem[p + 4] = arrayShift[3];
            if (NArea > 5) heapMem[p + 5] = arrayShift[4];
            if (NArea > 6) heapMem[p + 6] = arrayShift[5];
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          4: fork
            if (NArea > 4) heapMem[p + 4] = source1Value;
            if (NArea > 5) heapMem[p + 5] = arrayShift[4];
            if (NArea > 6) heapMem[p + 6] = arrayShift[5];
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          5: fork
            if (NArea > 5) heapMem[p + 5] = source1Value;
            if (NArea > 6) heapMem[p + 6] = arrayShift[5];
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          6: fork
            if (NArea > 6) heapMem[p + 6] = source1Value;
            if (NArea > 7) heapMem[p + 7] = arrayShift[6];
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          7: fork
            if (NArea > 7) heapMem[p + 7] = source1Value;
            if (NArea > 8) heapMem[p + 8] = arrayShift[7];
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          8: fork
            if (NArea > 8) heapMem[p + 8] = source1Value;
            if (NArea > 9) heapMem[p + 9] = arrayShift[8];
          join
          9: fork
            if (NArea > 9) heapMem[p + 9] = source1Value;
          join
        endcase
      end
    end
  endtask

  task moveLong_instruction();
    begin                                                                       // moveLong
      l = source2Value;
      p = targetLocation; j = sourceLocation;
      q = p + l;
      for(i = p; i < q; ++i) begin
        heapMem[i] = heapMem[j];
        ++j;
      end
    end
  endtask

  task in_instruction();
    begin                                                                       // in
     result = inMem[inMemPos++];
     setMemory();
    end
  endtask

  task inSize_instruction();
    begin                                                                       // inSize
     result = inMemEnd - inMemPos;
     setMemory();
    end
  endtask
endmodule
