//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire run,                                                              // Run - clock at lest once to allow code to be loaded
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  parameter integer MemoryElementWidth =  12;                                   // Memory element width

  parameter integer NArea   = 6;                                           // Size of each area on the heap
  parameter integer NArrays = 15;                                         // Maximum number of arrays
  parameter integer NHeap   = 6*15;                                  // Amount of heap memory
  parameter integer NLocal  = 2747;                                          // Size of local memory
  parameter integer NOut    =  2000;                                            // Size of output area
  parameter integer NIn            =     0;                                       // Size of input area
  reg [MemoryElementWidth-1:0]   arraySizes[NArrays-1:0];                       // Size of each array
  reg [MemoryElementWidth-1:0]      heapMem[NHeap-1  :0];                       // Heap memory
  reg [MemoryElementWidth-1:0]     localMem[NLocal-1 :0];                       // Local memory
  reg [MemoryElementWidth-1:0]       outMem[NOut-1   :0];                       // Out channel
  reg [MemoryElementWidth-1:0]        inMem[NIn-1    :0];                       // In channel
  reg [MemoryElementWidth-1:0]  freedArrays[NArrays-1:0];                       // Freed arrays list implemented as a stack
  reg [MemoryElementWidth-1:0]   arrayShift[NArea-1  :0];                       // Array shift area

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel
  integer allocs;                                                               // Maximum number of array allocations in use at any one time
  integer freedArraysTop;                                                       // Position in freed arrays stack

  integer ip;                                                                   // Instruction pointer
  reg     clock;                                                                // Clock - has to be one bit wide for yosys
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  task updateArrayLength(input integer arena, input integer array, input integer index); // Update array length if we are updating an array
    begin
      if (arena == 1 && arraySizes[array] < index + 1) arraySizes[array] = index + 1;
    end
  endtask

  always @(posedge run) begin                                                   // Initialize
    ip             = 0;
    clock          = 0;
    steps          = 0;
    finished       = 0;
    success        = 0;
    inMemPos       = 0;
    outMemPos      = 0;
    allocs         = 0;
    freedArraysTop = 0;
    for(i = 0; i < NHeap;   ++i)    heapMem[i] = 0;
    for(i = 0; i < NLocal;  ++i)   localMem[i] = 0;
    for(i = 0; i < NArrays; ++i) arraySizes[i] = 0;
  end

  always @(clock) begin                                                         // Each instruction
    steps = steps + 1;
    case(ip)

          0 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[0] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[0] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[0]] = 0;
              ip = 1;
      end

          1 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 2] = 3;
              updateArrayLength(1, localMem[0], 2);
              ip = 2;
      end

          2 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = 0;
              updateArrayLength(1, localMem[0], 3);
              ip = 3;
      end

          3 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = 0;
              updateArrayLength(1, localMem[0], 0);
              ip = 4;
      end

          4 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = 0;
              updateArrayLength(1, localMem[0], 1);
              ip = 5;
      end

          5 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1]] = 0;
              ip = 6;
      end

          6 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 7;
      end

          7 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 8;
      end

          8 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2] != 0 ? 31 : 9;
      end

          9 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[3] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[3] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[3]] = 0;
              ip = 10;
      end

         10 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 0] = 1;
              updateArrayLength(1, localMem[3], 0);
              ip = 11;
      end

         11 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 2] = 0;
              updateArrayLength(1, localMem[3], 2);
              ip = 12;
      end

         12 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[4] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[4] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[4]] = 0;
              ip = 13;
      end

         13 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 4] = localMem[4];
              updateArrayLength(1, localMem[3], 4);
              ip = 14;
      end

         14 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[5] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[5] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[5]] = 0;
              ip = 15;
      end

         15 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 5] = localMem[5];
              updateArrayLength(1, localMem[3], 5);
              ip = 16;
      end

         16 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 6] = 0;
              updateArrayLength(1, localMem[3], 6);
              ip = 17;
      end

         17 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 3] = localMem[0];
              updateArrayLength(1, localMem[3], 3);
              ip = 18;
      end

         18 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = heapMem[localMem[0]*6 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 19;
      end

         19 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*6 + 1] = heapMem[localMem[0]*6 + 1];
              updateArrayLength(1, localMem[3], 1);
              ip = 20;
      end

         20 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[6] = heapMem[localMem[3]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 21;
      end

         21 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[6]*6 + 0] = 1;
              updateArrayLength(1, localMem[6], 0);
              ip = 22;
      end

         22 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[7] = heapMem[localMem[3]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 23;
      end

         23 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[7]*6 + 0] = 11;
              updateArrayLength(1, localMem[7], 0);
              ip = 24;
      end

         24 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 25;
      end

         25 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = localMem[3];
              updateArrayLength(1, localMem[0], 3);
              ip = 26;
      end

         26 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[8] = heapMem[localMem[3]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 27;
      end

         27 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[8]] = 1;
              ip = 28;
      end

         28 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[9] = heapMem[localMem[3]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 29;
      end

         29 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[9]] = 1;
              ip = 30;
      end

         30 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1059;
      end

         31 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 32;
      end

         32 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[10] = heapMem[localMem[2]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 33;
      end

         33 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[11] = heapMem[localMem[0]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 34;
      end

         34 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[10] >= localMem[11] ? 70 : 35;
      end

         35 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[12] = heapMem[localMem[2]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 36;
      end

         36 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[12] != 0 ? 69 : 37;
      end

         37 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[13] = !heapMem[localMem[2]*6 + 6];
              ip = 38;
      end

         38 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[13] == 0 ? 68 : 39;
      end

         39 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[14] = heapMem[localMem[2]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 40;
      end

         40 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[15] = 0; k = arraySizes[localMem[14]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[14] * NArea + i] == 1) localMem[15] = i + 1;
              end
              ip = 41;
      end

         41 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[15] == 0 ? 46 : 42;
      end

         42 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[15] = localMem[15] - 1;
              updateArrayLength(2, 0, 0);
              ip = 43;
      end

         43 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[16] = heapMem[localMem[2]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 44;
      end

         44 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[16]*6 + localMem[15]] = 11;
              updateArrayLength(1, localMem[16], localMem[15]);
              ip = 45;
      end

         45 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1059;
      end

         46 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 47;
      end

         47 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[14]] = localMem[10];
              ip = 48;
      end

         48 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[17] = heapMem[localMem[2]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 49;
      end

         49 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[17]] = localMem[10];
              ip = 50;
      end

         50 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[14]];
//$display("AAAAA k=%d  source2=%d", k, 1);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[14] * NArea + i]);
                if (i < k && heapMem[localMem[14] * NArea + i] > 1) j = j + 1;
              end
              localMem[18] = j;
              ip = 51;
      end

         51 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[18] != 0 ? 59 : 52;
      end

         52 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[19] = heapMem[localMem[2]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 53;
      end

         53 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[19]*6 + localMem[10]] = 1;
              updateArrayLength(1, localMem[19], localMem[10]);
              ip = 54;
      end

         54 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[20] = heapMem[localMem[2]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 55;
      end

         55 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[20]*6 + localMem[10]] = 11;
              updateArrayLength(1, localMem[20], localMem[10]);
              ip = 56;
      end

         56 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2]*6 + 0] = localMem[10] + 1;
              updateArrayLength(1, localMem[2], 0);
              ip = 57;
      end

         57 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 58;
      end

         58 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1059;
      end

         59 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 60;
      end

         60 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[14]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[14] * NArea + i] < 1) j = j + 1;
              end
              localMem[21] = j;
              ip = 61;
      end

         61 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[22] = heapMem[localMem[2]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 62;
      end

         62 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[22] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[21], localMem[22], arraySizes[localMem[22]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[21] && i <= arraySizes[localMem[22]]) begin
                  heapMem[NArea * localMem[22] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[22] + localMem[21]] = 1;                                    // Insert new value
              arraySizes[localMem[22]] = arraySizes[localMem[22]] + 1;                              // Increase array size
              ip = 63;
      end

         63 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[23] = heapMem[localMem[2]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 64;
      end

         64 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[23] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[21], localMem[23], arraySizes[localMem[23]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[21] && i <= arraySizes[localMem[23]]) begin
                  heapMem[NArea * localMem[23] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[23] + localMem[21]] = 11;                                    // Insert new value
              arraySizes[localMem[23]] = arraySizes[localMem[23]] + 1;                              // Increase array size
              ip = 65;
      end

         65 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2]*6 + 0] = heapMem[localMem[2]*6 + 0] + 1;
              updateArrayLength(1, localMem[2], 0);
              ip = 66;
      end

         66 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 67;
      end

         67 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1059;
      end

         68 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 69;
      end

         69 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 70;
      end

         70 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 71;
      end

         71 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[24] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 72;
      end

         72 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 73;
      end

         73 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[26] = heapMem[localMem[24]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 74;
      end

         74 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[27] = heapMem[localMem[24]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 75;
      end

         75 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[28] = heapMem[localMem[27]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 76;
      end

         76 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[26] <  localMem[28] ? 296 : 77;
      end

         77 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[29] = localMem[28];
              updateArrayLength(2, 0, 0);
              ip = 78;
      end

         78 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[29] = localMem[29] >> 1;
              ip = 79;
      end

         79 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[30] = localMem[29] + 1;
              updateArrayLength(2, 0, 0);
              ip = 80;
      end

         80 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[31] = heapMem[localMem[24]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 81;
      end

         81 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[31] == 0 ? 178 : 82;
      end

         82 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[32] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[32] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[32]] = 0;
              ip = 83;
      end

         83 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 0] = localMem[29];
              updateArrayLength(1, localMem[32], 0);
              ip = 84;
      end

         84 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 2] = 0;
              updateArrayLength(1, localMem[32], 2);
              ip = 85;
      end

         85 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[33] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[33] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[33]] = 0;
              ip = 86;
      end

         86 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 4] = localMem[33];
              updateArrayLength(1, localMem[32], 4);
              ip = 87;
      end

         87 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[34] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[34] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[34]] = 0;
              ip = 88;
      end

         88 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 5] = localMem[34];
              updateArrayLength(1, localMem[32], 5);
              ip = 89;
      end

         89 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 6] = 0;
              updateArrayLength(1, localMem[32], 6);
              ip = 90;
      end

         90 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 3] = localMem[27];
              updateArrayLength(1, localMem[32], 3);
              ip = 91;
      end

         91 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[27]*6 + 1] = heapMem[localMem[27]*6 + 1] + 1;
              updateArrayLength(1, localMem[27], 1);
              ip = 92;
      end

         92 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 1] = heapMem[localMem[27]*6 + 1];
              updateArrayLength(1, localMem[32], 1);
              ip = 93;
      end

         93 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[35] = !heapMem[localMem[24]*6 + 6];
              ip = 94;
      end

         94 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[35] != 0 ? 123 : 95;
      end

         95 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[36] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[36] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[36]] = 0;
              ip = 96;
      end

         96 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 6] = localMem[36];
              updateArrayLength(1, localMem[32], 6);
              ip = 97;
      end

         97 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[37] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 98;
      end

         98 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[38] = heapMem[localMem[32]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 99;
      end

         99 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[38] + 0 + i] = heapMem[NArea * localMem[37] + localMem[30] + i];
                  updateArrayLength(1, localMem[38], 0 + i);
                end
              end
              ip = 100;
      end

        100 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[39] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 101;
      end

        101 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[40] = heapMem[localMem[32]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 102;
      end

        102 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[40] + 0 + i] = heapMem[NArea * localMem[39] + localMem[30] + i];
                  updateArrayLength(1, localMem[40], 0 + i);
                end
              end
              ip = 103;
      end

        103 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[41] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 104;
      end

        104 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[42] = heapMem[localMem[32]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 105;
      end

        105 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[43] = localMem[29] + 1;
              updateArrayLength(2, 0, 0);
              ip = 106;
      end

        106 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[43]) begin
                  heapMem[NArea * localMem[42] + 0 + i] = heapMem[NArea * localMem[41] + localMem[30] + i];
                  updateArrayLength(1, localMem[42], 0 + i);
                end
              end
              ip = 107;
      end

        107 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[44] = heapMem[localMem[32]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 108;
      end

        108 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[45] = localMem[44] + 1;
              updateArrayLength(2, 0, 0);
              ip = 109;
      end

        109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[46] = heapMem[localMem[32]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 110;
      end

        110 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 111;
      end

        111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[47] = 0;
              updateArrayLength(2, 0, 0);
              ip = 112;
      end

        112 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 113;
      end

        113 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[47] >= localMem[45] ? 119 : 114;
      end

        114 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[48] = heapMem[localMem[46]*6 + localMem[47]];
              updateArrayLength(2, 0, 0);
              ip = 115;
      end

        115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[48]*6 + 2] = localMem[32];
              updateArrayLength(1, localMem[48], 2);
              ip = 116;
      end

        116 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 117;
      end

        117 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[47] = localMem[47] + 1;
              updateArrayLength(2, 0, 0);
              ip = 118;
      end

        118 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 112;
      end

        119 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 120;
      end

        120 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[49] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 121;
      end

        121 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[49]] = localMem[30];
              ip = 122;
      end

        122 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 130;
      end

        123 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 124;
      end

        124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[50] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 125;
      end

        125 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[51] = heapMem[localMem[32]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 126;
      end

        126 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[51] + 0 + i] = heapMem[NArea * localMem[50] + localMem[30] + i];
                  updateArrayLength(1, localMem[51], 0 + i);
                end
              end
              ip = 127;
      end

        127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[52] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 128;
      end

        128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[53] = heapMem[localMem[32]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 129;
      end

        129 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[53] + 0 + i] = heapMem[NArea * localMem[52] + localMem[30] + i];
                  updateArrayLength(1, localMem[53], 0 + i);
                end
              end
              ip = 130;
      end

        130 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 131;
      end

        131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[24]*6 + 0] = localMem[29];
              updateArrayLength(1, localMem[24], 0);
              ip = 132;
      end

        132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[32]*6 + 2] = localMem[31];
              updateArrayLength(1, localMem[32], 2);
              ip = 133;
      end

        133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[54] = heapMem[localMem[31]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 134;
      end

        134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[55] = heapMem[localMem[31]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 135;
      end

        135 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[56] = heapMem[localMem[55]*6 + localMem[54]];
              updateArrayLength(2, 0, 0);
              ip = 136;
      end

        136 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[56] != localMem[24] ? 155 : 137;
      end

        137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[57] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 138;
      end

        138 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[58] = heapMem[localMem[57]*6 + localMem[29]];
              updateArrayLength(2, 0, 0);
              ip = 139;
      end

        139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[59] = heapMem[localMem[31]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 140;
      end

        140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[59]*6 + localMem[54]] = localMem[58];
              updateArrayLength(1, localMem[59], localMem[54]);
              ip = 141;
      end

        141 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[60] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 142;
      end

        142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[61] = heapMem[localMem[60]*6 + localMem[29]];
              updateArrayLength(2, 0, 0);
              ip = 143;
      end

        143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[62] = heapMem[localMem[31]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 144;
      end

        144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[62]*6 + localMem[54]] = localMem[61];
              updateArrayLength(1, localMem[62], localMem[54]);
              ip = 145;
      end

        145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[63] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 146;
      end

        146 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[63]] = localMem[29];
              ip = 147;
      end

        147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[64] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 148;
      end

        148 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[64]] = localMem[29];
              ip = 149;
      end

        149 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[65] = localMem[54] + 1;
              updateArrayLength(2, 0, 0);
              ip = 150;
      end

        150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[31]*6 + 0] = localMem[65];
              updateArrayLength(1, localMem[31], 0);
              ip = 151;
      end

        151 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[66] = heapMem[localMem[31]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 152;
      end

        152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[66]*6 + localMem[65]] = localMem[32];
              updateArrayLength(1, localMem[66], localMem[65]);
              ip = 153;
      end

        153 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 293;
      end

        154 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 177;
      end

        155 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 156;
      end

        156 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 157;
      end

        157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[67] = heapMem[localMem[31]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 158;
      end

        158 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[68] = 0; k = arraySizes[localMem[67]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[67] * NArea + i] == localMem[24]) localMem[68] = i + 1;
              end
              ip = 159;
      end

        159 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[68] = localMem[68] - 1;
              updateArrayLength(2, 0, 0);
              ip = 160;
      end

        160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[69] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 161;
      end

        161 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[70] = heapMem[localMem[69]*6 + localMem[29]];
              updateArrayLength(2, 0, 0);
              ip = 162;
      end

        162 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[71] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 163;
      end

        163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[72] = heapMem[localMem[71]*6 + localMem[29]];
              updateArrayLength(2, 0, 0);
              ip = 164;
      end

        164 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[73] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 165;
      end

        165 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[73]] = localMem[29];
              ip = 166;
      end

        166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[74] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 167;
      end

        167 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[74]] = localMem[29];
              ip = 168;
      end

        168 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[75] = heapMem[localMem[31]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 169;
      end

        169 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[75] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[68], localMem[75], arraySizes[localMem[75]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[68] && i <= arraySizes[localMem[75]]) begin
                  heapMem[NArea * localMem[75] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[75] + localMem[68]] = localMem[70];                                    // Insert new value
              arraySizes[localMem[75]] = arraySizes[localMem[75]] + 1;                              // Increase array size
              ip = 170;
      end

        170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[76] = heapMem[localMem[31]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 171;
      end

        171 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[76] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[68], localMem[76], arraySizes[localMem[76]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[68] && i <= arraySizes[localMem[76]]) begin
                  heapMem[NArea * localMem[76] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[76] + localMem[68]] = localMem[72];                                    // Insert new value
              arraySizes[localMem[76]] = arraySizes[localMem[76]] + 1;                              // Increase array size
              ip = 172;
      end

        172 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[77] = heapMem[localMem[31]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 173;
      end

        173 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[78] = localMem[68] + 1;
              updateArrayLength(2, 0, 0);
              ip = 174;
      end

        174 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[77] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[78], localMem[77], arraySizes[localMem[77]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[78] && i <= arraySizes[localMem[77]]) begin
                  heapMem[NArea * localMem[77] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[77] + localMem[78]] = localMem[32];                                    // Insert new value
              arraySizes[localMem[77]] = arraySizes[localMem[77]] + 1;                              // Increase array size
              ip = 175;
      end

        175 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[31]*6 + 0] = heapMem[localMem[31]*6 + 0] + 1;
              updateArrayLength(1, localMem[31], 0);
              ip = 176;
      end

        176 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 293;
      end

        177 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 178;
      end

        178 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 179;
      end

        179 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[79] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[79] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[79]] = 0;
              ip = 180;
      end

        180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 0] = localMem[29];
              updateArrayLength(1, localMem[79], 0);
              ip = 181;
      end

        181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 2] = 0;
              updateArrayLength(1, localMem[79], 2);
              ip = 182;
      end

        182 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[80] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[80] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[80]] = 0;
              ip = 183;
      end

        183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 4] = localMem[80];
              updateArrayLength(1, localMem[79], 4);
              ip = 184;
      end

        184 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[81] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[81] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[81]] = 0;
              ip = 185;
      end

        185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 5] = localMem[81];
              updateArrayLength(1, localMem[79], 5);
              ip = 186;
      end

        186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 6] = 0;
              updateArrayLength(1, localMem[79], 6);
              ip = 187;
      end

        187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 3] = localMem[27];
              updateArrayLength(1, localMem[79], 3);
              ip = 188;
      end

        188 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[27]*6 + 1] = heapMem[localMem[27]*6 + 1] + 1;
              updateArrayLength(1, localMem[27], 1);
              ip = 189;
      end

        189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 1] = heapMem[localMem[27]*6 + 1];
              updateArrayLength(1, localMem[79], 1);
              ip = 190;
      end

        190 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[82] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[82] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[82]] = 0;
              ip = 191;
      end

        191 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 0] = localMem[29];
              updateArrayLength(1, localMem[82], 0);
              ip = 192;
      end

        192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 2] = 0;
              updateArrayLength(1, localMem[82], 2);
              ip = 193;
      end

        193 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[83] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[83] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[83]] = 0;
              ip = 194;
      end

        194 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 4] = localMem[83];
              updateArrayLength(1, localMem[82], 4);
              ip = 195;
      end

        195 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[84] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[84] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[84]] = 0;
              ip = 196;
      end

        196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 5] = localMem[84];
              updateArrayLength(1, localMem[82], 5);
              ip = 197;
      end

        197 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 6] = 0;
              updateArrayLength(1, localMem[82], 6);
              ip = 198;
      end

        198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 3] = localMem[27];
              updateArrayLength(1, localMem[82], 3);
              ip = 199;
      end

        199 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[27]*6 + 1] = heapMem[localMem[27]*6 + 1] + 1;
              updateArrayLength(1, localMem[27], 1);
              ip = 200;
      end

        200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 1] = heapMem[localMem[27]*6 + 1];
              updateArrayLength(1, localMem[82], 1);
              ip = 201;
      end

        201 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[85] = !heapMem[localMem[24]*6 + 6];
              ip = 202;
      end

        202 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[85] != 0 ? 254 : 203;
      end

        203 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[86] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[86] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[86]] = 0;
              ip = 204;
      end

        204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 6] = localMem[86];
              updateArrayLength(1, localMem[79], 6);
              ip = 205;
      end

        205 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[87] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[87] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[87]] = 0;
              ip = 206;
      end

        206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 6] = localMem[87];
              updateArrayLength(1, localMem[82], 6);
              ip = 207;
      end

        207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[88] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 208;
      end

        208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[89] = heapMem[localMem[79]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 209;
      end

        209 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[89] + 0 + i] = heapMem[NArea * localMem[88] + 0 + i];
                  updateArrayLength(1, localMem[89], 0 + i);
                end
              end
              ip = 210;
      end

        210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[90] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 211;
      end

        211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[91] = heapMem[localMem[79]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 212;
      end

        212 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[91] + 0 + i] = heapMem[NArea * localMem[90] + 0 + i];
                  updateArrayLength(1, localMem[91], 0 + i);
                end
              end
              ip = 213;
      end

        213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[92] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 214;
      end

        214 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[93] = heapMem[localMem[79]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 215;
      end

        215 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[94] = localMem[29] + 1;
              updateArrayLength(2, 0, 0);
              ip = 216;
      end

        216 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[94]) begin
                  heapMem[NArea * localMem[93] + 0 + i] = heapMem[NArea * localMem[92] + 0 + i];
                  updateArrayLength(1, localMem[93], 0 + i);
                end
              end
              ip = 217;
      end

        217 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[95] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 218;
      end

        218 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[96] = heapMem[localMem[82]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 219;
      end

        219 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[96] + 0 + i] = heapMem[NArea * localMem[95] + localMem[30] + i];
                  updateArrayLength(1, localMem[96], 0 + i);
                end
              end
              ip = 220;
      end

        220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[97] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 221;
      end

        221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[98] = heapMem[localMem[82]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 222;
      end

        222 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[98] + 0 + i] = heapMem[NArea * localMem[97] + localMem[30] + i];
                  updateArrayLength(1, localMem[98], 0 + i);
                end
              end
              ip = 223;
      end

        223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[99] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 224;
      end

        224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[100] = heapMem[localMem[82]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 225;
      end

        225 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[101] = localMem[29] + 1;
              updateArrayLength(2, 0, 0);
              ip = 226;
      end

        226 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[101]) begin
                  heapMem[NArea * localMem[100] + 0 + i] = heapMem[NArea * localMem[99] + localMem[30] + i];
                  updateArrayLength(1, localMem[100], 0 + i);
                end
              end
              ip = 227;
      end

        227 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[102] = heapMem[localMem[79]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 228;
      end

        228 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[103] = localMem[102] + 1;
              updateArrayLength(2, 0, 0);
              ip = 229;
      end

        229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[104] = heapMem[localMem[79]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 230;
      end

        230 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 231;
      end

        231 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[105] = 0;
              updateArrayLength(2, 0, 0);
              ip = 232;
      end

        232 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 233;
      end

        233 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[105] >= localMem[103] ? 239 : 234;
      end

        234 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[106] = heapMem[localMem[104]*6 + localMem[105]];
              updateArrayLength(2, 0, 0);
              ip = 235;
      end

        235 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[106]*6 + 2] = localMem[79];
              updateArrayLength(1, localMem[106], 2);
              ip = 236;
      end

        236 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 237;
      end

        237 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[105] = localMem[105] + 1;
              updateArrayLength(2, 0, 0);
              ip = 238;
      end

        238 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 232;
      end

        239 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 240;
      end

        240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[107] = heapMem[localMem[82]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 241;
      end

        241 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[108] = localMem[107] + 1;
              updateArrayLength(2, 0, 0);
              ip = 242;
      end

        242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[109] = heapMem[localMem[82]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 243;
      end

        243 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 244;
      end

        244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[110] = 0;
              updateArrayLength(2, 0, 0);
              ip = 245;
      end

        245 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 246;
      end

        246 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[110] >= localMem[108] ? 252 : 247;
      end

        247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[111] = heapMem[localMem[109]*6 + localMem[110]];
              updateArrayLength(2, 0, 0);
              ip = 248;
      end

        248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[111]*6 + 2] = localMem[82];
              updateArrayLength(1, localMem[111], 2);
              ip = 249;
      end

        249 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 250;
      end

        250 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[110] = localMem[110] + 1;
              updateArrayLength(2, 0, 0);
              ip = 251;
      end

        251 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 245;
      end

        252 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 253;
      end

        253 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 269;
      end

        254 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 255;
      end

        255 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[112] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[112] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[112]] = 0;
              ip = 256;
      end

        256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[24]*6 + 6] = localMem[112];
              updateArrayLength(1, localMem[24], 6);
              ip = 257;
      end

        257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[113] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 258;
      end

        258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[114] = heapMem[localMem[79]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 259;
      end

        259 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[114] + 0 + i] = heapMem[NArea * localMem[113] + 0 + i];
                  updateArrayLength(1, localMem[114], 0 + i);
                end
              end
              ip = 260;
      end

        260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[115] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 261;
      end

        261 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[116] = heapMem[localMem[79]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 262;
      end

        262 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[116] + 0 + i] = heapMem[NArea * localMem[115] + 0 + i];
                  updateArrayLength(1, localMem[116], 0 + i);
                end
              end
              ip = 263;
      end

        263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[117] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 264;
      end

        264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[118] = heapMem[localMem[82]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 265;
      end

        265 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[118] + 0 + i] = heapMem[NArea * localMem[117] + localMem[30] + i];
                  updateArrayLength(1, localMem[118], 0 + i);
                end
              end
              ip = 266;
      end

        266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[119] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 267;
      end

        267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[120] = heapMem[localMem[82]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 268;
      end

        268 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[29]) begin
                  heapMem[NArea * localMem[120] + 0 + i] = heapMem[NArea * localMem[119] + localMem[30] + i];
                  updateArrayLength(1, localMem[120], 0 + i);
                end
              end
              ip = 269;
      end

        269 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 270;
      end

        270 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[79]*6 + 2] = localMem[24];
              updateArrayLength(1, localMem[79], 2);
              ip = 271;
      end

        271 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[82]*6 + 2] = localMem[24];
              updateArrayLength(1, localMem[82], 2);
              ip = 272;
      end

        272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[121] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 273;
      end

        273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[122] = heapMem[localMem[121]*6 + localMem[29]];
              updateArrayLength(2, 0, 0);
              ip = 274;
      end

        274 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[123] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 275;
      end

        275 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[124] = heapMem[localMem[123]*6 + localMem[29]];
              updateArrayLength(2, 0, 0);
              ip = 276;
      end

        276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[125] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 277;
      end

        277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[125]*6 + 0] = localMem[122];
              updateArrayLength(1, localMem[125], 0);
              ip = 278;
      end

        278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[126] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 279;
      end

        279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[126]*6 + 0] = localMem[124];
              updateArrayLength(1, localMem[126], 0);
              ip = 280;
      end

        280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[127] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 281;
      end

        281 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[127]*6 + 0] = localMem[79];
              updateArrayLength(1, localMem[127], 0);
              ip = 282;
      end

        282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[128] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 283;
      end

        283 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[128]*6 + 1] = localMem[82];
              updateArrayLength(1, localMem[128], 1);
              ip = 284;
      end

        284 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[24]*6 + 0] = 1;
              updateArrayLength(1, localMem[24], 0);
              ip = 285;
      end

        285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[129] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 286;
      end

        286 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[129]] = 1;
              ip = 287;
      end

        287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[130] = heapMem[localMem[24]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 288;
      end

        288 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[130]] = 1;
              ip = 289;
      end

        289 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[131] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 290;
      end

        290 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[131]] = 2;
              ip = 291;
      end

        291 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 293;
      end

        292 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 298;
      end

        293 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 294;
      end

        294 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[25] = 1;
              updateArrayLength(2, 0, 0);
              ip = 295;
      end

        295 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 298;
      end

        296 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 297;
      end

        297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[25] = 0;
              updateArrayLength(2, 0, 0);
              ip = 298;
      end

        298 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 299;
      end

        299 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 300;
      end

        300 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 301;
      end

        301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[132] = 0;
              updateArrayLength(2, 0, 0);
              ip = 302;
      end

        302 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 303;
      end

        303 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[132] >= 99 ? 801 : 304;
      end

        304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[133] = heapMem[localMem[24]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 305;
      end

        305 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[134] = localMem[133] - 1;
              updateArrayLength(2, 0, 0);
              ip = 306;
      end

        306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[135] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 307;
      end

        307 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[136] = heapMem[localMem[135]*6 + localMem[134]];
              updateArrayLength(2, 0, 0);
              ip = 308;
      end

        308 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 1 <= localMem[136] ? 549 : 309;
      end

        309 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[137] = !heapMem[localMem[24]*6 + 6];
              ip = 310;
      end

        310 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[137] == 0 ? 315 : 311;
      end

        311 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 0] = localMem[24];
              updateArrayLength(1, localMem[1], 0);
              ip = 312;
      end

        312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 1] = 2;
              updateArrayLength(1, localMem[1], 1);
              ip = 313;
      end

        313 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1]*6 + 2] = localMem[133] - 1;
              updateArrayLength(1, localMem[1], 2);
              ip = 314;
      end

        314 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 805;
      end

        315 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 316;
      end

        316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[138] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 317;
      end

        317 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[139] = heapMem[localMem[138]*6 + localMem[133]];
              updateArrayLength(2, 0, 0);
              ip = 318;
      end

        318 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 319;
      end

        319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[141] = heapMem[localMem[139]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 320;
      end

        320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[142] = heapMem[localMem[139]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 321;
      end

        321 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[143] = heapMem[localMem[142]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 322;
      end

        322 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[141] <  localMem[143] ? 542 : 323;
      end

        323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[144] = localMem[143];
              updateArrayLength(2, 0, 0);
              ip = 324;
      end

        324 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[144] = localMem[144] >> 1;
              ip = 325;
      end

        325 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[145] = localMem[144] + 1;
              updateArrayLength(2, 0, 0);
              ip = 326;
      end

        326 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[146] = heapMem[localMem[139]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 327;
      end

        327 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[146] == 0 ? 424 : 328;
      end

        328 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[147] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[147] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[147]] = 0;
              ip = 329;
      end

        329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 0] = localMem[144];
              updateArrayLength(1, localMem[147], 0);
              ip = 330;
      end

        330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 2] = 0;
              updateArrayLength(1, localMem[147], 2);
              ip = 331;
      end

        331 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[148] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[148] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[148]] = 0;
              ip = 332;
      end

        332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 4] = localMem[148];
              updateArrayLength(1, localMem[147], 4);
              ip = 333;
      end

        333 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[149] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[149] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[149]] = 0;
              ip = 334;
      end

        334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 5] = localMem[149];
              updateArrayLength(1, localMem[147], 5);
              ip = 335;
      end

        335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 6] = 0;
              updateArrayLength(1, localMem[147], 6);
              ip = 336;
      end

        336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 3] = localMem[142];
              updateArrayLength(1, localMem[147], 3);
              ip = 337;
      end

        337 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[142]*6 + 1] = heapMem[localMem[142]*6 + 1] + 1;
              updateArrayLength(1, localMem[142], 1);
              ip = 338;
      end

        338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 1] = heapMem[localMem[142]*6 + 1];
              updateArrayLength(1, localMem[147], 1);
              ip = 339;
      end

        339 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[150] = !heapMem[localMem[139]*6 + 6];
              ip = 340;
      end

        340 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[150] != 0 ? 369 : 341;
      end

        341 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[151] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[151] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[151]] = 0;
              ip = 342;
      end

        342 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 6] = localMem[151];
              updateArrayLength(1, localMem[147], 6);
              ip = 343;
      end

        343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[152] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 344;
      end

        344 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[153] = heapMem[localMem[147]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 345;
      end

        345 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[153] + 0 + i] = heapMem[NArea * localMem[152] + localMem[145] + i];
                  updateArrayLength(1, localMem[153], 0 + i);
                end
              end
              ip = 346;
      end

        346 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[154] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 347;
      end

        347 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[155] = heapMem[localMem[147]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 348;
      end

        348 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[155] + 0 + i] = heapMem[NArea * localMem[154] + localMem[145] + i];
                  updateArrayLength(1, localMem[155], 0 + i);
                end
              end
              ip = 349;
      end

        349 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[156] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 350;
      end

        350 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[157] = heapMem[localMem[147]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 351;
      end

        351 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[158] = localMem[144] + 1;
              updateArrayLength(2, 0, 0);
              ip = 352;
      end

        352 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[158]) begin
                  heapMem[NArea * localMem[157] + 0 + i] = heapMem[NArea * localMem[156] + localMem[145] + i];
                  updateArrayLength(1, localMem[157], 0 + i);
                end
              end
              ip = 353;
      end

        353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[159] = heapMem[localMem[147]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 354;
      end

        354 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[160] = localMem[159] + 1;
              updateArrayLength(2, 0, 0);
              ip = 355;
      end

        355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[161] = heapMem[localMem[147]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 356;
      end

        356 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 357;
      end

        357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[162] = 0;
              updateArrayLength(2, 0, 0);
              ip = 358;
      end

        358 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 359;
      end

        359 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[162] >= localMem[160] ? 365 : 360;
      end

        360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[163] = heapMem[localMem[161]*6 + localMem[162]];
              updateArrayLength(2, 0, 0);
              ip = 361;
      end

        361 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[163]*6 + 2] = localMem[147];
              updateArrayLength(1, localMem[163], 2);
              ip = 362;
      end

        362 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 363;
      end

        363 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[162] = localMem[162] + 1;
              updateArrayLength(2, 0, 0);
              ip = 364;
      end

        364 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 358;
      end

        365 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 366;
      end

        366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[164] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 367;
      end

        367 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[164]] = localMem[145];
              ip = 368;
      end

        368 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 376;
      end

        369 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 370;
      end

        370 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[165] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 371;
      end

        371 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[166] = heapMem[localMem[147]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 372;
      end

        372 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[166] + 0 + i] = heapMem[NArea * localMem[165] + localMem[145] + i];
                  updateArrayLength(1, localMem[166], 0 + i);
                end
              end
              ip = 373;
      end

        373 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[167] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 374;
      end

        374 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[168] = heapMem[localMem[147]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 375;
      end

        375 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[168] + 0 + i] = heapMem[NArea * localMem[167] + localMem[145] + i];
                  updateArrayLength(1, localMem[168], 0 + i);
                end
              end
              ip = 376;
      end

        376 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 377;
      end

        377 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[139]*6 + 0] = localMem[144];
              updateArrayLength(1, localMem[139], 0);
              ip = 378;
      end

        378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[147]*6 + 2] = localMem[146];
              updateArrayLength(1, localMem[147], 2);
              ip = 379;
      end

        379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[169] = heapMem[localMem[146]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 380;
      end

        380 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[170] = heapMem[localMem[146]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 381;
      end

        381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[171] = heapMem[localMem[170]*6 + localMem[169]];
              updateArrayLength(2, 0, 0);
              ip = 382;
      end

        382 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[171] != localMem[139] ? 401 : 383;
      end

        383 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[172] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 384;
      end

        384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[173] = heapMem[localMem[172]*6 + localMem[144]];
              updateArrayLength(2, 0, 0);
              ip = 385;
      end

        385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[174] = heapMem[localMem[146]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 386;
      end

        386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[174]*6 + localMem[169]] = localMem[173];
              updateArrayLength(1, localMem[174], localMem[169]);
              ip = 387;
      end

        387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[175] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 388;
      end

        388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[176] = heapMem[localMem[175]*6 + localMem[144]];
              updateArrayLength(2, 0, 0);
              ip = 389;
      end

        389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[177] = heapMem[localMem[146]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 390;
      end

        390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[177]*6 + localMem[169]] = localMem[176];
              updateArrayLength(1, localMem[177], localMem[169]);
              ip = 391;
      end

        391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[178] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 392;
      end

        392 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[178]] = localMem[144];
              ip = 393;
      end

        393 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[179] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 394;
      end

        394 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[179]] = localMem[144];
              ip = 395;
      end

        395 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[180] = localMem[169] + 1;
              updateArrayLength(2, 0, 0);
              ip = 396;
      end

        396 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[146]*6 + 0] = localMem[180];
              updateArrayLength(1, localMem[146], 0);
              ip = 397;
      end

        397 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[181] = heapMem[localMem[146]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 398;
      end

        398 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[181]*6 + localMem[180]] = localMem[147];
              updateArrayLength(1, localMem[181], localMem[180]);
              ip = 399;
      end

        399 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 539;
      end

        400 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 423;
      end

        401 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 402;
      end

        402 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 403;
      end

        403 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[182] = heapMem[localMem[146]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 404;
      end

        404 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[183] = 0; k = arraySizes[localMem[182]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[182] * NArea + i] == localMem[139]) localMem[183] = i + 1;
              end
              ip = 405;
      end

        405 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[183] = localMem[183] - 1;
              updateArrayLength(2, 0, 0);
              ip = 406;
      end

        406 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[184] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 407;
      end

        407 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[185] = heapMem[localMem[184]*6 + localMem[144]];
              updateArrayLength(2, 0, 0);
              ip = 408;
      end

        408 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[186] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 409;
      end

        409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[187] = heapMem[localMem[186]*6 + localMem[144]];
              updateArrayLength(2, 0, 0);
              ip = 410;
      end

        410 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[188] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 411;
      end

        411 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[188]] = localMem[144];
              ip = 412;
      end

        412 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[189] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 413;
      end

        413 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[189]] = localMem[144];
              ip = 414;
      end

        414 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[190] = heapMem[localMem[146]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 415;
      end

        415 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[190] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[183], localMem[190], arraySizes[localMem[190]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[183] && i <= arraySizes[localMem[190]]) begin
                  heapMem[NArea * localMem[190] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[190] + localMem[183]] = localMem[185];                                    // Insert new value
              arraySizes[localMem[190]] = arraySizes[localMem[190]] + 1;                              // Increase array size
              ip = 416;
      end

        416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[191] = heapMem[localMem[146]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 417;
      end

        417 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[191] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[183], localMem[191], arraySizes[localMem[191]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[183] && i <= arraySizes[localMem[191]]) begin
                  heapMem[NArea * localMem[191] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[191] + localMem[183]] = localMem[187];                                    // Insert new value
              arraySizes[localMem[191]] = arraySizes[localMem[191]] + 1;                              // Increase array size
              ip = 418;
      end

        418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[192] = heapMem[localMem[146]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 419;
      end

        419 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[193] = localMem[183] + 1;
              updateArrayLength(2, 0, 0);
              ip = 420;
      end

        420 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[192] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[193], localMem[192], arraySizes[localMem[192]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[193] && i <= arraySizes[localMem[192]]) begin
                  heapMem[NArea * localMem[192] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[192] + localMem[193]] = localMem[147];                                    // Insert new value
              arraySizes[localMem[192]] = arraySizes[localMem[192]] + 1;                              // Increase array size
              ip = 421;
      end

        421 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[146]*6 + 0] = heapMem[localMem[146]*6 + 0] + 1;
              updateArrayLength(1, localMem[146], 0);
              ip = 422;
      end

        422 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 539;
      end

        423 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 424;
      end

        424 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 425;
      end

        425 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[194] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[194] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[194]] = 0;
              ip = 426;
      end

        426 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 0] = localMem[144];
              updateArrayLength(1, localMem[194], 0);
              ip = 427;
      end

        427 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 2] = 0;
              updateArrayLength(1, localMem[194], 2);
              ip = 428;
      end

        428 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[195] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[195] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[195]] = 0;
              ip = 429;
      end

        429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 4] = localMem[195];
              updateArrayLength(1, localMem[194], 4);
              ip = 430;
      end

        430 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[196] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[196] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[196]] = 0;
              ip = 431;
      end

        431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 5] = localMem[196];
              updateArrayLength(1, localMem[194], 5);
              ip = 432;
      end

        432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 6] = 0;
              updateArrayLength(1, localMem[194], 6);
              ip = 433;
      end

        433 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 3] = localMem[142];
              updateArrayLength(1, localMem[194], 3);
              ip = 434;
      end

        434 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[142]*6 + 1] = heapMem[localMem[142]*6 + 1] + 1;
              updateArrayLength(1, localMem[142], 1);
              ip = 435;
      end

        435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 1] = heapMem[localMem[142]*6 + 1];
              updateArrayLength(1, localMem[194], 1);
              ip = 436;
      end

        436 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[197] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[197] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[197]] = 0;
              ip = 437;
      end

        437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 0] = localMem[144];
              updateArrayLength(1, localMem[197], 0);
              ip = 438;
      end

        438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 2] = 0;
              updateArrayLength(1, localMem[197], 2);
              ip = 439;
      end

        439 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[198] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[198] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[198]] = 0;
              ip = 440;
      end

        440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 4] = localMem[198];
              updateArrayLength(1, localMem[197], 4);
              ip = 441;
      end

        441 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[199] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[199] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[199]] = 0;
              ip = 442;
      end

        442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 5] = localMem[199];
              updateArrayLength(1, localMem[197], 5);
              ip = 443;
      end

        443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 6] = 0;
              updateArrayLength(1, localMem[197], 6);
              ip = 444;
      end

        444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 3] = localMem[142];
              updateArrayLength(1, localMem[197], 3);
              ip = 445;
      end

        445 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[142]*6 + 1] = heapMem[localMem[142]*6 + 1] + 1;
              updateArrayLength(1, localMem[142], 1);
              ip = 446;
      end

        446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 1] = heapMem[localMem[142]*6 + 1];
              updateArrayLength(1, localMem[197], 1);
              ip = 447;
      end

        447 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[200] = !heapMem[localMem[139]*6 + 6];
              ip = 448;
      end

        448 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[200] != 0 ? 500 : 449;
      end

        449 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[201] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[201] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[201]] = 0;
              ip = 450;
      end

        450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 6] = localMem[201];
              updateArrayLength(1, localMem[194], 6);
              ip = 451;
      end

        451 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[202] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[202] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[202]] = 0;
              ip = 452;
      end

        452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 6] = localMem[202];
              updateArrayLength(1, localMem[197], 6);
              ip = 453;
      end

        453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[203] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 454;
      end

        454 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[204] = heapMem[localMem[194]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 455;
      end

        455 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[204] + 0 + i] = heapMem[NArea * localMem[203] + 0 + i];
                  updateArrayLength(1, localMem[204], 0 + i);
                end
              end
              ip = 456;
      end

        456 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[205] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 457;
      end

        457 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[206] = heapMem[localMem[194]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 458;
      end

        458 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[206] + 0 + i] = heapMem[NArea * localMem[205] + 0 + i];
                  updateArrayLength(1, localMem[206], 0 + i);
                end
              end
              ip = 459;
      end

        459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[207] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 460;
      end

        460 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[208] = heapMem[localMem[194]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 461;
      end

        461 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[209] = localMem[144] + 1;
              updateArrayLength(2, 0, 0);
              ip = 462;
      end

        462 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[209]) begin
                  heapMem[NArea * localMem[208] + 0 + i] = heapMem[NArea * localMem[207] + 0 + i];
                  updateArrayLength(1, localMem[208], 0 + i);
                end
              end
              ip = 463;
      end

        463 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[210] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 464;
      end

        464 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[211] = heapMem[localMem[197]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 465;
      end

        465 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[211] + 0 + i] = heapMem[NArea * localMem[210] + localMem[145] + i];
                  updateArrayLength(1, localMem[211], 0 + i);
                end
              end
              ip = 466;
      end

        466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[212] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 467;
      end

        467 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[213] = heapMem[localMem[197]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 468;
      end

        468 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[213] + 0 + i] = heapMem[NArea * localMem[212] + localMem[145] + i];
                  updateArrayLength(1, localMem[213], 0 + i);
                end
              end
              ip = 469;
      end

        469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[214] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 470;
      end

        470 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[215] = heapMem[localMem[197]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 471;
      end

        471 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[216] = localMem[144] + 1;
              updateArrayLength(2, 0, 0);
              ip = 472;
      end

        472 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[216]) begin
                  heapMem[NArea * localMem[215] + 0 + i] = heapMem[NArea * localMem[214] + localMem[145] + i];
                  updateArrayLength(1, localMem[215], 0 + i);
                end
              end
              ip = 473;
      end

        473 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[217] = heapMem[localMem[194]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 474;
      end

        474 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[218] = localMem[217] + 1;
              updateArrayLength(2, 0, 0);
              ip = 475;
      end

        475 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[219] = heapMem[localMem[194]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 476;
      end

        476 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 477;
      end

        477 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[220] = 0;
              updateArrayLength(2, 0, 0);
              ip = 478;
      end

        478 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 479;
      end

        479 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[220] >= localMem[218] ? 485 : 480;
      end

        480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[221] = heapMem[localMem[219]*6 + localMem[220]];
              updateArrayLength(2, 0, 0);
              ip = 481;
      end

        481 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[221]*6 + 2] = localMem[194];
              updateArrayLength(1, localMem[221], 2);
              ip = 482;
      end

        482 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 483;
      end

        483 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[220] = localMem[220] + 1;
              updateArrayLength(2, 0, 0);
              ip = 484;
      end

        484 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 478;
      end

        485 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 486;
      end

        486 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[222] = heapMem[localMem[197]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 487;
      end

        487 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[223] = localMem[222] + 1;
              updateArrayLength(2, 0, 0);
              ip = 488;
      end

        488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[224] = heapMem[localMem[197]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 489;
      end

        489 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 490;
      end

        490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[225] = 0;
              updateArrayLength(2, 0, 0);
              ip = 491;
      end

        491 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 492;
      end

        492 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[225] >= localMem[223] ? 498 : 493;
      end

        493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[226] = heapMem[localMem[224]*6 + localMem[225]];
              updateArrayLength(2, 0, 0);
              ip = 494;
      end

        494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[226]*6 + 2] = localMem[197];
              updateArrayLength(1, localMem[226], 2);
              ip = 495;
      end

        495 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 496;
      end

        496 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[225] = localMem[225] + 1;
              updateArrayLength(2, 0, 0);
              ip = 497;
      end

        497 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 491;
      end

        498 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 499;
      end

        499 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 515;
      end

        500 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 501;
      end

        501 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[227] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[227] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[227]] = 0;
              ip = 502;
      end

        502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[139]*6 + 6] = localMem[227];
              updateArrayLength(1, localMem[139], 6);
              ip = 503;
      end

        503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[228] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 504;
      end

        504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[229] = heapMem[localMem[194]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 505;
      end

        505 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[229] + 0 + i] = heapMem[NArea * localMem[228] + 0 + i];
                  updateArrayLength(1, localMem[229], 0 + i);
                end
              end
              ip = 506;
      end

        506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[230] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 507;
      end

        507 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[231] = heapMem[localMem[194]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 508;
      end

        508 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[231] + 0 + i] = heapMem[NArea * localMem[230] + 0 + i];
                  updateArrayLength(1, localMem[231], 0 + i);
                end
              end
              ip = 509;
      end

        509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[232] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 510;
      end

        510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[233] = heapMem[localMem[197]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 511;
      end

        511 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[233] + 0 + i] = heapMem[NArea * localMem[232] + localMem[145] + i];
                  updateArrayLength(1, localMem[233], 0 + i);
                end
              end
              ip = 512;
      end

        512 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[234] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 513;
      end

        513 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[235] = heapMem[localMem[197]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 514;
      end

        514 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[144]) begin
                  heapMem[NArea * localMem[235] + 0 + i] = heapMem[NArea * localMem[234] + localMem[145] + i];
                  updateArrayLength(1, localMem[235], 0 + i);
                end
              end
              ip = 515;
      end

        515 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 516;
      end

        516 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[194]*6 + 2] = localMem[139];
              updateArrayLength(1, localMem[194], 2);
              ip = 517;
      end

        517 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[197]*6 + 2] = localMem[139];
              updateArrayLength(1, localMem[197], 2);
              ip = 518;
      end

        518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[236] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 519;
      end

        519 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[237] = heapMem[localMem[236]*6 + localMem[144]];
              updateArrayLength(2, 0, 0);
              ip = 520;
      end

        520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[238] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 521;
      end

        521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[239] = heapMem[localMem[238]*6 + localMem[144]];
              updateArrayLength(2, 0, 0);
              ip = 522;
      end

        522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[240] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 523;
      end

        523 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[240]*6 + 0] = localMem[237];
              updateArrayLength(1, localMem[240], 0);
              ip = 524;
      end

        524 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[241] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 525;
      end

        525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[241]*6 + 0] = localMem[239];
              updateArrayLength(1, localMem[241], 0);
              ip = 526;
      end

        526 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[242] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 527;
      end

        527 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[242]*6 + 0] = localMem[194];
              updateArrayLength(1, localMem[242], 0);
              ip = 528;
      end

        528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[243] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 529;
      end

        529 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[243]*6 + 1] = localMem[197];
              updateArrayLength(1, localMem[243], 1);
              ip = 530;
      end

        530 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[139]*6 + 0] = 1;
              updateArrayLength(1, localMem[139], 0);
              ip = 531;
      end

        531 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[244] = heapMem[localMem[139]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 532;
      end

        532 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[244]] = 1;
              ip = 533;
      end

        533 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[245] = heapMem[localMem[139]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 534;
      end

        534 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[245]] = 1;
              ip = 535;
      end

        535 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[246] = heapMem[localMem[139]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 536;
      end

        536 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[246]] = 2;
              ip = 537;
      end

        537 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 539;
      end

        538 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 544;
      end

        539 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 540;
      end

        540 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[140] = 1;
              updateArrayLength(2, 0, 0);
              ip = 541;
      end

        541 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 544;
      end

        542 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 543;
      end

        543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[140] = 0;
              updateArrayLength(2, 0, 0);
              ip = 544;
      end

        544 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 545;
      end

        545 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[140] != 0 ? 547 : 546;
      end

        546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[24] = localMem[139];
              updateArrayLength(2, 0, 0);
              ip = 547;
      end

        547 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 548;
      end

        548 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 798;
      end

        549 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 550;
      end

        550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[247] = heapMem[localMem[24]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 551;
      end

        551 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[248] = 0; k = arraySizes[localMem[247]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[247] * NArea + i] == 1) localMem[248] = i + 1;
              end
              ip = 552;
      end

        552 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[248] == 0 ? 557 : 553;
      end

        553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 0] = localMem[24];
              updateArrayLength(1, localMem[1], 0);
              ip = 554;
      end

        554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 1] = 1;
              updateArrayLength(1, localMem[1], 1);
              ip = 555;
      end

        555 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1]*6 + 2] = localMem[248] - 1;
              updateArrayLength(1, localMem[1], 2);
              ip = 556;
      end

        556 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 805;
      end

        557 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 558;
      end

        558 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[247]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[247] * NArea + i] < 1) j = j + 1;
              end
              localMem[249] = j;
              ip = 559;
      end

        559 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[250] = !heapMem[localMem[24]*6 + 6];
              ip = 560;
      end

        560 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[250] == 0 ? 565 : 561;
      end

        561 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 0] = localMem[24];
              updateArrayLength(1, localMem[1], 0);
              ip = 562;
      end

        562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 1] = 0;
              updateArrayLength(1, localMem[1], 1);
              ip = 563;
      end

        563 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1]*6 + 2] = localMem[249];
              updateArrayLength(1, localMem[1], 2);
              ip = 564;
      end

        564 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 805;
      end

        565 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 566;
      end

        566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[251] = heapMem[localMem[24]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 567;
      end

        567 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[252] = heapMem[localMem[251]*6 + localMem[249]];
              updateArrayLength(2, 0, 0);
              ip = 568;
      end

        568 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 569;
      end

        569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[254] = heapMem[localMem[252]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 570;
      end

        570 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[255] = heapMem[localMem[252]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 571;
      end

        571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[256] = heapMem[localMem[255]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 572;
      end

        572 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[254] <  localMem[256] ? 792 : 573;
      end

        573 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[257] = localMem[256];
              updateArrayLength(2, 0, 0);
              ip = 574;
      end

        574 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[257] = localMem[257] >> 1;
              ip = 575;
      end

        575 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[258] = localMem[257] + 1;
              updateArrayLength(2, 0, 0);
              ip = 576;
      end

        576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[259] = heapMem[localMem[252]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 577;
      end

        577 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[259] == 0 ? 674 : 578;
      end

        578 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[260] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[260] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[260]] = 0;
              ip = 579;
      end

        579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 0] = localMem[257];
              updateArrayLength(1, localMem[260], 0);
              ip = 580;
      end

        580 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 2] = 0;
              updateArrayLength(1, localMem[260], 2);
              ip = 581;
      end

        581 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[261] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[261] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[261]] = 0;
              ip = 582;
      end

        582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 4] = localMem[261];
              updateArrayLength(1, localMem[260], 4);
              ip = 583;
      end

        583 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[262] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[262] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[262]] = 0;
              ip = 584;
      end

        584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 5] = localMem[262];
              updateArrayLength(1, localMem[260], 5);
              ip = 585;
      end

        585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 6] = 0;
              updateArrayLength(1, localMem[260], 6);
              ip = 586;
      end

        586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 3] = localMem[255];
              updateArrayLength(1, localMem[260], 3);
              ip = 587;
      end

        587 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[255]*6 + 1] = heapMem[localMem[255]*6 + 1] + 1;
              updateArrayLength(1, localMem[255], 1);
              ip = 588;
      end

        588 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 1] = heapMem[localMem[255]*6 + 1];
              updateArrayLength(1, localMem[260], 1);
              ip = 589;
      end

        589 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[263] = !heapMem[localMem[252]*6 + 6];
              ip = 590;
      end

        590 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[263] != 0 ? 619 : 591;
      end

        591 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[264] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[264] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[264]] = 0;
              ip = 592;
      end

        592 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 6] = localMem[264];
              updateArrayLength(1, localMem[260], 6);
              ip = 593;
      end

        593 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[265] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 594;
      end

        594 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[266] = heapMem[localMem[260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 595;
      end

        595 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[266] + 0 + i] = heapMem[NArea * localMem[265] + localMem[258] + i];
                  updateArrayLength(1, localMem[266], 0 + i);
                end
              end
              ip = 596;
      end

        596 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[267] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 597;
      end

        597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[268] = heapMem[localMem[260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 598;
      end

        598 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[268] + 0 + i] = heapMem[NArea * localMem[267] + localMem[258] + i];
                  updateArrayLength(1, localMem[268], 0 + i);
                end
              end
              ip = 599;
      end

        599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[269] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 600;
      end

        600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[270] = heapMem[localMem[260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 601;
      end

        601 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[271] = localMem[257] + 1;
              updateArrayLength(2, 0, 0);
              ip = 602;
      end

        602 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[271]) begin
                  heapMem[NArea * localMem[270] + 0 + i] = heapMem[NArea * localMem[269] + localMem[258] + i];
                  updateArrayLength(1, localMem[270], 0 + i);
                end
              end
              ip = 603;
      end

        603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[272] = heapMem[localMem[260]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 604;
      end

        604 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[273] = localMem[272] + 1;
              updateArrayLength(2, 0, 0);
              ip = 605;
      end

        605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[274] = heapMem[localMem[260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 606;
      end

        606 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 607;
      end

        607 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[275] = 0;
              updateArrayLength(2, 0, 0);
              ip = 608;
      end

        608 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 609;
      end

        609 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[275] >= localMem[273] ? 615 : 610;
      end

        610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[276] = heapMem[localMem[274]*6 + localMem[275]];
              updateArrayLength(2, 0, 0);
              ip = 611;
      end

        611 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[276]*6 + 2] = localMem[260];
              updateArrayLength(1, localMem[276], 2);
              ip = 612;
      end

        612 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 613;
      end

        613 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[275] = localMem[275] + 1;
              updateArrayLength(2, 0, 0);
              ip = 614;
      end

        614 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 608;
      end

        615 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 616;
      end

        616 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[277] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 617;
      end

        617 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[277]] = localMem[258];
              ip = 618;
      end

        618 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 626;
      end

        619 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 620;
      end

        620 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[278] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 621;
      end

        621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[279] = heapMem[localMem[260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 622;
      end

        622 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[279] + 0 + i] = heapMem[NArea * localMem[278] + localMem[258] + i];
                  updateArrayLength(1, localMem[279], 0 + i);
                end
              end
              ip = 623;
      end

        623 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[280] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 624;
      end

        624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[281] = heapMem[localMem[260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 625;
      end

        625 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[281] + 0 + i] = heapMem[NArea * localMem[280] + localMem[258] + i];
                  updateArrayLength(1, localMem[281], 0 + i);
                end
              end
              ip = 626;
      end

        626 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 627;
      end

        627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[252]*6 + 0] = localMem[257];
              updateArrayLength(1, localMem[252], 0);
              ip = 628;
      end

        628 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[260]*6 + 2] = localMem[259];
              updateArrayLength(1, localMem[260], 2);
              ip = 629;
      end

        629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[282] = heapMem[localMem[259]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 630;
      end

        630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[283] = heapMem[localMem[259]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 631;
      end

        631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[284] = heapMem[localMem[283]*6 + localMem[282]];
              updateArrayLength(2, 0, 0);
              ip = 632;
      end

        632 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[284] != localMem[252] ? 651 : 633;
      end

        633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[285] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 634;
      end

        634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[286] = heapMem[localMem[285]*6 + localMem[257]];
              updateArrayLength(2, 0, 0);
              ip = 635;
      end

        635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[287] = heapMem[localMem[259]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 636;
      end

        636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[287]*6 + localMem[282]] = localMem[286];
              updateArrayLength(1, localMem[287], localMem[282]);
              ip = 637;
      end

        637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[288] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 638;
      end

        638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[289] = heapMem[localMem[288]*6 + localMem[257]];
              updateArrayLength(2, 0, 0);
              ip = 639;
      end

        639 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[290] = heapMem[localMem[259]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 640;
      end

        640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[290]*6 + localMem[282]] = localMem[289];
              updateArrayLength(1, localMem[290], localMem[282]);
              ip = 641;
      end

        641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[291] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 642;
      end

        642 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[291]] = localMem[257];
              ip = 643;
      end

        643 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[292] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 644;
      end

        644 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[292]] = localMem[257];
              ip = 645;
      end

        645 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[293] = localMem[282] + 1;
              updateArrayLength(2, 0, 0);
              ip = 646;
      end

        646 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[259]*6 + 0] = localMem[293];
              updateArrayLength(1, localMem[259], 0);
              ip = 647;
      end

        647 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[294] = heapMem[localMem[259]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 648;
      end

        648 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[294]*6 + localMem[293]] = localMem[260];
              updateArrayLength(1, localMem[294], localMem[293]);
              ip = 649;
      end

        649 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 789;
      end

        650 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 673;
      end

        651 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 652;
      end

        652 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 653;
      end

        653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[295] = heapMem[localMem[259]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 654;
      end

        654 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[296] = 0; k = arraySizes[localMem[295]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[295] * NArea + i] == localMem[252]) localMem[296] = i + 1;
              end
              ip = 655;
      end

        655 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[296] = localMem[296] - 1;
              updateArrayLength(2, 0, 0);
              ip = 656;
      end

        656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[297] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 657;
      end

        657 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[298] = heapMem[localMem[297]*6 + localMem[257]];
              updateArrayLength(2, 0, 0);
              ip = 658;
      end

        658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[299] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 659;
      end

        659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[300] = heapMem[localMem[299]*6 + localMem[257]];
              updateArrayLength(2, 0, 0);
              ip = 660;
      end

        660 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[301] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 661;
      end

        661 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[301]] = localMem[257];
              ip = 662;
      end

        662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[302] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 663;
      end

        663 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[302]] = localMem[257];
              ip = 664;
      end

        664 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[303] = heapMem[localMem[259]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 665;
      end

        665 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[303] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[296], localMem[303], arraySizes[localMem[303]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[296] && i <= arraySizes[localMem[303]]) begin
                  heapMem[NArea * localMem[303] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[303] + localMem[296]] = localMem[298];                                    // Insert new value
              arraySizes[localMem[303]] = arraySizes[localMem[303]] + 1;                              // Increase array size
              ip = 666;
      end

        666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[304] = heapMem[localMem[259]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 667;
      end

        667 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[304] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[296], localMem[304], arraySizes[localMem[304]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[296] && i <= arraySizes[localMem[304]]) begin
                  heapMem[NArea * localMem[304] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[304] + localMem[296]] = localMem[300];                                    // Insert new value
              arraySizes[localMem[304]] = arraySizes[localMem[304]] + 1;                              // Increase array size
              ip = 668;
      end

        668 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[305] = heapMem[localMem[259]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 669;
      end

        669 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[306] = localMem[296] + 1;
              updateArrayLength(2, 0, 0);
              ip = 670;
      end

        670 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[305] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[306], localMem[305], arraySizes[localMem[305]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[306] && i <= arraySizes[localMem[305]]) begin
                  heapMem[NArea * localMem[305] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[305] + localMem[306]] = localMem[260];                                    // Insert new value
              arraySizes[localMem[305]] = arraySizes[localMem[305]] + 1;                              // Increase array size
              ip = 671;
      end

        671 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[259]*6 + 0] = heapMem[localMem[259]*6 + 0] + 1;
              updateArrayLength(1, localMem[259], 0);
              ip = 672;
      end

        672 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 789;
      end

        673 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 674;
      end

        674 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 675;
      end

        675 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[307] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[307] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[307]] = 0;
              ip = 676;
      end

        676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 0] = localMem[257];
              updateArrayLength(1, localMem[307], 0);
              ip = 677;
      end

        677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 2] = 0;
              updateArrayLength(1, localMem[307], 2);
              ip = 678;
      end

        678 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[308] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[308] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[308]] = 0;
              ip = 679;
      end

        679 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 4] = localMem[308];
              updateArrayLength(1, localMem[307], 4);
              ip = 680;
      end

        680 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[309] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[309] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[309]] = 0;
              ip = 681;
      end

        681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 5] = localMem[309];
              updateArrayLength(1, localMem[307], 5);
              ip = 682;
      end

        682 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 6] = 0;
              updateArrayLength(1, localMem[307], 6);
              ip = 683;
      end

        683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 3] = localMem[255];
              updateArrayLength(1, localMem[307], 3);
              ip = 684;
      end

        684 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[255]*6 + 1] = heapMem[localMem[255]*6 + 1] + 1;
              updateArrayLength(1, localMem[255], 1);
              ip = 685;
      end

        685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 1] = heapMem[localMem[255]*6 + 1];
              updateArrayLength(1, localMem[307], 1);
              ip = 686;
      end

        686 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[310] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[310] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[310]] = 0;
              ip = 687;
      end

        687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 0] = localMem[257];
              updateArrayLength(1, localMem[310], 0);
              ip = 688;
      end

        688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 2] = 0;
              updateArrayLength(1, localMem[310], 2);
              ip = 689;
      end

        689 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[311] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[311] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[311]] = 0;
              ip = 690;
      end

        690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 4] = localMem[311];
              updateArrayLength(1, localMem[310], 4);
              ip = 691;
      end

        691 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[312] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[312] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[312]] = 0;
              ip = 692;
      end

        692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 5] = localMem[312];
              updateArrayLength(1, localMem[310], 5);
              ip = 693;
      end

        693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 6] = 0;
              updateArrayLength(1, localMem[310], 6);
              ip = 694;
      end

        694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 3] = localMem[255];
              updateArrayLength(1, localMem[310], 3);
              ip = 695;
      end

        695 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[255]*6 + 1] = heapMem[localMem[255]*6 + 1] + 1;
              updateArrayLength(1, localMem[255], 1);
              ip = 696;
      end

        696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 1] = heapMem[localMem[255]*6 + 1];
              updateArrayLength(1, localMem[310], 1);
              ip = 697;
      end

        697 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[313] = !heapMem[localMem[252]*6 + 6];
              ip = 698;
      end

        698 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[313] != 0 ? 750 : 699;
      end

        699 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[314] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[314] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[314]] = 0;
              ip = 700;
      end

        700 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 6] = localMem[314];
              updateArrayLength(1, localMem[307], 6);
              ip = 701;
      end

        701 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[315] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[315] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[315]] = 0;
              ip = 702;
      end

        702 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 6] = localMem[315];
              updateArrayLength(1, localMem[310], 6);
              ip = 703;
      end

        703 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[316] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 704;
      end

        704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[317] = heapMem[localMem[307]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 705;
      end

        705 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[317] + 0 + i] = heapMem[NArea * localMem[316] + 0 + i];
                  updateArrayLength(1, localMem[317], 0 + i);
                end
              end
              ip = 706;
      end

        706 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[318] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 707;
      end

        707 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[319] = heapMem[localMem[307]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 708;
      end

        708 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[319] + 0 + i] = heapMem[NArea * localMem[318] + 0 + i];
                  updateArrayLength(1, localMem[319], 0 + i);
                end
              end
              ip = 709;
      end

        709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[320] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 710;
      end

        710 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[321] = heapMem[localMem[307]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 711;
      end

        711 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[322] = localMem[257] + 1;
              updateArrayLength(2, 0, 0);
              ip = 712;
      end

        712 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[322]) begin
                  heapMem[NArea * localMem[321] + 0 + i] = heapMem[NArea * localMem[320] + 0 + i];
                  updateArrayLength(1, localMem[321], 0 + i);
                end
              end
              ip = 713;
      end

        713 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[323] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 714;
      end

        714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[324] = heapMem[localMem[310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 715;
      end

        715 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[324] + 0 + i] = heapMem[NArea * localMem[323] + localMem[258] + i];
                  updateArrayLength(1, localMem[324], 0 + i);
                end
              end
              ip = 716;
      end

        716 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[325] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 717;
      end

        717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[326] = heapMem[localMem[310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 718;
      end

        718 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[326] + 0 + i] = heapMem[NArea * localMem[325] + localMem[258] + i];
                  updateArrayLength(1, localMem[326], 0 + i);
                end
              end
              ip = 719;
      end

        719 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[327] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 720;
      end

        720 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[328] = heapMem[localMem[310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 721;
      end

        721 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[329] = localMem[257] + 1;
              updateArrayLength(2, 0, 0);
              ip = 722;
      end

        722 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[329]) begin
                  heapMem[NArea * localMem[328] + 0 + i] = heapMem[NArea * localMem[327] + localMem[258] + i];
                  updateArrayLength(1, localMem[328], 0 + i);
                end
              end
              ip = 723;
      end

        723 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[330] = heapMem[localMem[307]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 724;
      end

        724 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[331] = localMem[330] + 1;
              updateArrayLength(2, 0, 0);
              ip = 725;
      end

        725 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[332] = heapMem[localMem[307]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 726;
      end

        726 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 727;
      end

        727 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[333] = 0;
              updateArrayLength(2, 0, 0);
              ip = 728;
      end

        728 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 729;
      end

        729 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[333] >= localMem[331] ? 735 : 730;
      end

        730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[334] = heapMem[localMem[332]*6 + localMem[333]];
              updateArrayLength(2, 0, 0);
              ip = 731;
      end

        731 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[334]*6 + 2] = localMem[307];
              updateArrayLength(1, localMem[334], 2);
              ip = 732;
      end

        732 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 733;
      end

        733 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[333] = localMem[333] + 1;
              updateArrayLength(2, 0, 0);
              ip = 734;
      end

        734 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 728;
      end

        735 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 736;
      end

        736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[335] = heapMem[localMem[310]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 737;
      end

        737 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[336] = localMem[335] + 1;
              updateArrayLength(2, 0, 0);
              ip = 738;
      end

        738 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[337] = heapMem[localMem[310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 739;
      end

        739 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 740;
      end

        740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[338] = 0;
              updateArrayLength(2, 0, 0);
              ip = 741;
      end

        741 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 742;
      end

        742 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[338] >= localMem[336] ? 748 : 743;
      end

        743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[339] = heapMem[localMem[337]*6 + localMem[338]];
              updateArrayLength(2, 0, 0);
              ip = 744;
      end

        744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[339]*6 + 2] = localMem[310];
              updateArrayLength(1, localMem[339], 2);
              ip = 745;
      end

        745 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 746;
      end

        746 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[338] = localMem[338] + 1;
              updateArrayLength(2, 0, 0);
              ip = 747;
      end

        747 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 741;
      end

        748 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 749;
      end

        749 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 765;
      end

        750 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 751;
      end

        751 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[340] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[340] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[340]] = 0;
              ip = 752;
      end

        752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[252]*6 + 6] = localMem[340];
              updateArrayLength(1, localMem[252], 6);
              ip = 753;
      end

        753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[341] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 754;
      end

        754 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[342] = heapMem[localMem[307]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 755;
      end

        755 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[342] + 0 + i] = heapMem[NArea * localMem[341] + 0 + i];
                  updateArrayLength(1, localMem[342], 0 + i);
                end
              end
              ip = 756;
      end

        756 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[343] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 757;
      end

        757 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[344] = heapMem[localMem[307]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 758;
      end

        758 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[344] + 0 + i] = heapMem[NArea * localMem[343] + 0 + i];
                  updateArrayLength(1, localMem[344], 0 + i);
                end
              end
              ip = 759;
      end

        759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[345] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 760;
      end

        760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[346] = heapMem[localMem[310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 761;
      end

        761 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[346] + 0 + i] = heapMem[NArea * localMem[345] + localMem[258] + i];
                  updateArrayLength(1, localMem[346], 0 + i);
                end
              end
              ip = 762;
      end

        762 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[347] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 763;
      end

        763 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[348] = heapMem[localMem[310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 764;
      end

        764 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[257]) begin
                  heapMem[NArea * localMem[348] + 0 + i] = heapMem[NArea * localMem[347] + localMem[258] + i];
                  updateArrayLength(1, localMem[348], 0 + i);
                end
              end
              ip = 765;
      end

        765 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 766;
      end

        766 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[307]*6 + 2] = localMem[252];
              updateArrayLength(1, localMem[307], 2);
              ip = 767;
      end

        767 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[310]*6 + 2] = localMem[252];
              updateArrayLength(1, localMem[310], 2);
              ip = 768;
      end

        768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[349] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 769;
      end

        769 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[350] = heapMem[localMem[349]*6 + localMem[257]];
              updateArrayLength(2, 0, 0);
              ip = 770;
      end

        770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[351] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 771;
      end

        771 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[352] = heapMem[localMem[351]*6 + localMem[257]];
              updateArrayLength(2, 0, 0);
              ip = 772;
      end

        772 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[353] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 773;
      end

        773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[353]*6 + 0] = localMem[350];
              updateArrayLength(1, localMem[353], 0);
              ip = 774;
      end

        774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[354] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 775;
      end

        775 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[354]*6 + 0] = localMem[352];
              updateArrayLength(1, localMem[354], 0);
              ip = 776;
      end

        776 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[355] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 777;
      end

        777 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[355]*6 + 0] = localMem[307];
              updateArrayLength(1, localMem[355], 0);
              ip = 778;
      end

        778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[356] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 779;
      end

        779 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[356]*6 + 1] = localMem[310];
              updateArrayLength(1, localMem[356], 1);
              ip = 780;
      end

        780 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[252]*6 + 0] = 1;
              updateArrayLength(1, localMem[252], 0);
              ip = 781;
      end

        781 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[357] = heapMem[localMem[252]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 782;
      end

        782 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[357]] = 1;
              ip = 783;
      end

        783 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[358] = heapMem[localMem[252]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 784;
      end

        784 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[358]] = 1;
              ip = 785;
      end

        785 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[359] = heapMem[localMem[252]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 786;
      end

        786 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[359]] = 2;
              ip = 787;
      end

        787 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 789;
      end

        788 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 794;
      end

        789 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 790;
      end

        790 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[253] = 1;
              updateArrayLength(2, 0, 0);
              ip = 791;
      end

        791 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 794;
      end

        792 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 793;
      end

        793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[253] = 0;
              updateArrayLength(2, 0, 0);
              ip = 794;
      end

        794 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 795;
      end

        795 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[253] != 0 ? 797 : 796;
      end

        796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[24] = localMem[252];
              updateArrayLength(2, 0, 0);
              ip = 797;
      end

        797 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 798;
      end

        798 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 799;
      end

        799 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[132] = localMem[132] + 1;
              updateArrayLength(2, 0, 0);
              ip = 800;
      end

        800 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 302;
      end

        801 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 802;
      end

        802 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
            ip = 803;
      end

        803 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 804;
      end

        804 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 805;
      end

        805 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 806;
      end

        806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[360] = heapMem[localMem[1]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 807;
      end

        807 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[361] = heapMem[localMem[1]*6 + 1];
              updateArrayLength(2, 0, 0);
              ip = 808;
      end

        808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[362] = heapMem[localMem[1]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 809;
      end

        809 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[361] != 1 ? 813 : 810;
      end

        810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[363] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 811;
      end

        811 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[363]*6 + localMem[362]] = 11;
              updateArrayLength(1, localMem[363], localMem[362]);
              ip = 812;
      end

        812 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1059;
      end

        813 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 814;
      end

        814 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[361] != 2 ? 822 : 815;
      end

        815 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[364] = localMem[362] + 1;
              updateArrayLength(2, 0, 0);
              ip = 816;
      end

        816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[365] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 817;
      end

        817 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[365] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[364], localMem[365], arraySizes[localMem[365]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[364] && i <= arraySizes[localMem[365]]) begin
                  heapMem[NArea * localMem[365] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[365] + localMem[364]] = 1;                                    // Insert new value
              arraySizes[localMem[365]] = arraySizes[localMem[365]] + 1;                              // Increase array size
              ip = 818;
      end

        818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[366] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 819;
      end

        819 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[366] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[364], localMem[366], arraySizes[localMem[366]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[364] && i <= arraySizes[localMem[366]]) begin
                  heapMem[NArea * localMem[366] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[366] + localMem[364]] = 11;                                    // Insert new value
              arraySizes[localMem[366]] = arraySizes[localMem[366]] + 1;                              // Increase array size
              ip = 820;
      end

        820 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[360]*6 + 0] = heapMem[localMem[360]*6 + 0] + 1;
              updateArrayLength(1, localMem[360], 0);
              ip = 821;
      end

        821 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 828;
      end

        822 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 823;
      end

        823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[367] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 824;
      end

        824 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[367] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[362], localMem[367], arraySizes[localMem[367]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[362] && i <= arraySizes[localMem[367]]) begin
                  heapMem[NArea * localMem[367] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[367] + localMem[362]] = 1;                                    // Insert new value
              arraySizes[localMem[367]] = arraySizes[localMem[367]] + 1;                              // Increase array size
              ip = 825;
      end

        825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[368] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 826;
      end

        826 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[368] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[362], localMem[368], arraySizes[localMem[368]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[362] && i <= arraySizes[localMem[368]]) begin
                  heapMem[NArea * localMem[368] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[368] + localMem[362]] = 11;                                    // Insert new value
              arraySizes[localMem[368]] = arraySizes[localMem[368]] + 1;                              // Increase array size
              ip = 827;
      end

        827 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[360]*6 + 0] = heapMem[localMem[360]*6 + 0] + 1;
              updateArrayLength(1, localMem[360], 0);
              ip = 828;
      end

        828 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 829;
      end

        829 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 830;
      end

        830 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 831;
      end

        831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[370] = heapMem[localMem[360]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 832;
      end

        832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[371] = heapMem[localMem[360]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 833;
      end

        833 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[372] = heapMem[localMem[371]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 834;
      end

        834 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[370] <  localMem[372] ? 1054 : 835;
      end

        835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[373] = localMem[372];
              updateArrayLength(2, 0, 0);
              ip = 836;
      end

        836 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[373] = localMem[373] >> 1;
              ip = 837;
      end

        837 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[374] = localMem[373] + 1;
              updateArrayLength(2, 0, 0);
              ip = 838;
      end

        838 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[375] = heapMem[localMem[360]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 839;
      end

        839 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[375] == 0 ? 936 : 840;
      end

        840 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[376] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[376] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[376]] = 0;
              ip = 841;
      end

        841 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 0] = localMem[373];
              updateArrayLength(1, localMem[376], 0);
              ip = 842;
      end

        842 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 2] = 0;
              updateArrayLength(1, localMem[376], 2);
              ip = 843;
      end

        843 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[377] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[377] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[377]] = 0;
              ip = 844;
      end

        844 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 4] = localMem[377];
              updateArrayLength(1, localMem[376], 4);
              ip = 845;
      end

        845 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[378] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[378] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[378]] = 0;
              ip = 846;
      end

        846 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 5] = localMem[378];
              updateArrayLength(1, localMem[376], 5);
              ip = 847;
      end

        847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 6] = 0;
              updateArrayLength(1, localMem[376], 6);
              ip = 848;
      end

        848 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 3] = localMem[371];
              updateArrayLength(1, localMem[376], 3);
              ip = 849;
      end

        849 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[371]*6 + 1] = heapMem[localMem[371]*6 + 1] + 1;
              updateArrayLength(1, localMem[371], 1);
              ip = 850;
      end

        850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 1] = heapMem[localMem[371]*6 + 1];
              updateArrayLength(1, localMem[376], 1);
              ip = 851;
      end

        851 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[379] = !heapMem[localMem[360]*6 + 6];
              ip = 852;
      end

        852 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[379] != 0 ? 881 : 853;
      end

        853 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[380] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[380] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[380]] = 0;
              ip = 854;
      end

        854 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 6] = localMem[380];
              updateArrayLength(1, localMem[376], 6);
              ip = 855;
      end

        855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[381] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 856;
      end

        856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[382] = heapMem[localMem[376]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 857;
      end

        857 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[382] + 0 + i] = heapMem[NArea * localMem[381] + localMem[374] + i];
                  updateArrayLength(1, localMem[382], 0 + i);
                end
              end
              ip = 858;
      end

        858 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[383] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 859;
      end

        859 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[384] = heapMem[localMem[376]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 860;
      end

        860 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[384] + 0 + i] = heapMem[NArea * localMem[383] + localMem[374] + i];
                  updateArrayLength(1, localMem[384], 0 + i);
                end
              end
              ip = 861;
      end

        861 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[385] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 862;
      end

        862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[386] = heapMem[localMem[376]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 863;
      end

        863 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[387] = localMem[373] + 1;
              updateArrayLength(2, 0, 0);
              ip = 864;
      end

        864 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[387]) begin
                  heapMem[NArea * localMem[386] + 0 + i] = heapMem[NArea * localMem[385] + localMem[374] + i];
                  updateArrayLength(1, localMem[386], 0 + i);
                end
              end
              ip = 865;
      end

        865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[388] = heapMem[localMem[376]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 866;
      end

        866 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[389] = localMem[388] + 1;
              updateArrayLength(2, 0, 0);
              ip = 867;
      end

        867 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[390] = heapMem[localMem[376]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 868;
      end

        868 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 869;
      end

        869 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[391] = 0;
              updateArrayLength(2, 0, 0);
              ip = 870;
      end

        870 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 871;
      end

        871 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[391] >= localMem[389] ? 877 : 872;
      end

        872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[392] = heapMem[localMem[390]*6 + localMem[391]];
              updateArrayLength(2, 0, 0);
              ip = 873;
      end

        873 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[392]*6 + 2] = localMem[376];
              updateArrayLength(1, localMem[392], 2);
              ip = 874;
      end

        874 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 875;
      end

        875 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[391] = localMem[391] + 1;
              updateArrayLength(2, 0, 0);
              ip = 876;
      end

        876 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 870;
      end

        877 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 878;
      end

        878 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[393] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 879;
      end

        879 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[393]] = localMem[374];
              ip = 880;
      end

        880 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 888;
      end

        881 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 882;
      end

        882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[394] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 883;
      end

        883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[395] = heapMem[localMem[376]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 884;
      end

        884 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[395] + 0 + i] = heapMem[NArea * localMem[394] + localMem[374] + i];
                  updateArrayLength(1, localMem[395], 0 + i);
                end
              end
              ip = 885;
      end

        885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[396] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 886;
      end

        886 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[397] = heapMem[localMem[376]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 887;
      end

        887 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[397] + 0 + i] = heapMem[NArea * localMem[396] + localMem[374] + i];
                  updateArrayLength(1, localMem[397], 0 + i);
                end
              end
              ip = 888;
      end

        888 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 889;
      end

        889 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[360]*6 + 0] = localMem[373];
              updateArrayLength(1, localMem[360], 0);
              ip = 890;
      end

        890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[376]*6 + 2] = localMem[375];
              updateArrayLength(1, localMem[376], 2);
              ip = 891;
      end

        891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[398] = heapMem[localMem[375]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 892;
      end

        892 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[399] = heapMem[localMem[375]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 893;
      end

        893 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[400] = heapMem[localMem[399]*6 + localMem[398]];
              updateArrayLength(2, 0, 0);
              ip = 894;
      end

        894 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[400] != localMem[360] ? 913 : 895;
      end

        895 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[401] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 896;
      end

        896 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[402] = heapMem[localMem[401]*6 + localMem[373]];
              updateArrayLength(2, 0, 0);
              ip = 897;
      end

        897 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[403] = heapMem[localMem[375]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 898;
      end

        898 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[403]*6 + localMem[398]] = localMem[402];
              updateArrayLength(1, localMem[403], localMem[398]);
              ip = 899;
      end

        899 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[404] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 900;
      end

        900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[405] = heapMem[localMem[404]*6 + localMem[373]];
              updateArrayLength(2, 0, 0);
              ip = 901;
      end

        901 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[406] = heapMem[localMem[375]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 902;
      end

        902 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[406]*6 + localMem[398]] = localMem[405];
              updateArrayLength(1, localMem[406], localMem[398]);
              ip = 903;
      end

        903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[407] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 904;
      end

        904 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[407]] = localMem[373];
              ip = 905;
      end

        905 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[408] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 906;
      end

        906 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[408]] = localMem[373];
              ip = 907;
      end

        907 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[409] = localMem[398] + 1;
              updateArrayLength(2, 0, 0);
              ip = 908;
      end

        908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[375]*6 + 0] = localMem[409];
              updateArrayLength(1, localMem[375], 0);
              ip = 909;
      end

        909 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[410] = heapMem[localMem[375]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 910;
      end

        910 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[410]*6 + localMem[409]] = localMem[376];
              updateArrayLength(1, localMem[410], localMem[409]);
              ip = 911;
      end

        911 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1051;
      end

        912 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 935;
      end

        913 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 914;
      end

        914 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 915;
      end

        915 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[411] = heapMem[localMem[375]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 916;
      end

        916 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[412] = 0; k = arraySizes[localMem[411]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[411] * NArea + i] == localMem[360]) localMem[412] = i + 1;
              end
              ip = 917;
      end

        917 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[412] = localMem[412] - 1;
              updateArrayLength(2, 0, 0);
              ip = 918;
      end

        918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[413] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 919;
      end

        919 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[414] = heapMem[localMem[413]*6 + localMem[373]];
              updateArrayLength(2, 0, 0);
              ip = 920;
      end

        920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[415] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 921;
      end

        921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[416] = heapMem[localMem[415]*6 + localMem[373]];
              updateArrayLength(2, 0, 0);
              ip = 922;
      end

        922 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[417] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 923;
      end

        923 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[417]] = localMem[373];
              ip = 924;
      end

        924 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[418] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 925;
      end

        925 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[418]] = localMem[373];
              ip = 926;
      end

        926 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[419] = heapMem[localMem[375]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 927;
      end

        927 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[419] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[412], localMem[419], arraySizes[localMem[419]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[412] && i <= arraySizes[localMem[419]]) begin
                  heapMem[NArea * localMem[419] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[419] + localMem[412]] = localMem[414];                                    // Insert new value
              arraySizes[localMem[419]] = arraySizes[localMem[419]] + 1;                              // Increase array size
              ip = 928;
      end

        928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[420] = heapMem[localMem[375]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 929;
      end

        929 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[420] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[412], localMem[420], arraySizes[localMem[420]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[412] && i <= arraySizes[localMem[420]]) begin
                  heapMem[NArea * localMem[420] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[420] + localMem[412]] = localMem[416];                                    // Insert new value
              arraySizes[localMem[420]] = arraySizes[localMem[420]] + 1;                              // Increase array size
              ip = 930;
      end

        930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[421] = heapMem[localMem[375]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 931;
      end

        931 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[422] = localMem[412] + 1;
              updateArrayLength(2, 0, 0);
              ip = 932;
      end

        932 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[421] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[422], localMem[421], arraySizes[localMem[421]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[422] && i <= arraySizes[localMem[421]]) begin
                  heapMem[NArea * localMem[421] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[421] + localMem[422]] = localMem[376];                                    // Insert new value
              arraySizes[localMem[421]] = arraySizes[localMem[421]] + 1;                              // Increase array size
              ip = 933;
      end

        933 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[375]*6 + 0] = heapMem[localMem[375]*6 + 0] + 1;
              updateArrayLength(1, localMem[375], 0);
              ip = 934;
      end

        934 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1051;
      end

        935 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 936;
      end

        936 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 937;
      end

        937 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[423] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[423] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[423]] = 0;
              ip = 938;
      end

        938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 0] = localMem[373];
              updateArrayLength(1, localMem[423], 0);
              ip = 939;
      end

        939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 2] = 0;
              updateArrayLength(1, localMem[423], 2);
              ip = 940;
      end

        940 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[424] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[424] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[424]] = 0;
              ip = 941;
      end

        941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 4] = localMem[424];
              updateArrayLength(1, localMem[423], 4);
              ip = 942;
      end

        942 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[425] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[425] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[425]] = 0;
              ip = 943;
      end

        943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 5] = localMem[425];
              updateArrayLength(1, localMem[423], 5);
              ip = 944;
      end

        944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 6] = 0;
              updateArrayLength(1, localMem[423], 6);
              ip = 945;
      end

        945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 3] = localMem[371];
              updateArrayLength(1, localMem[423], 3);
              ip = 946;
      end

        946 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[371]*6 + 1] = heapMem[localMem[371]*6 + 1] + 1;
              updateArrayLength(1, localMem[371], 1);
              ip = 947;
      end

        947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 1] = heapMem[localMem[371]*6 + 1];
              updateArrayLength(1, localMem[423], 1);
              ip = 948;
      end

        948 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[426] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[426] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[426]] = 0;
              ip = 949;
      end

        949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 0] = localMem[373];
              updateArrayLength(1, localMem[426], 0);
              ip = 950;
      end

        950 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 2] = 0;
              updateArrayLength(1, localMem[426], 2);
              ip = 951;
      end

        951 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[427] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[427] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[427]] = 0;
              ip = 952;
      end

        952 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 4] = localMem[427];
              updateArrayLength(1, localMem[426], 4);
              ip = 953;
      end

        953 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[428] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[428] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[428]] = 0;
              ip = 954;
      end

        954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 5] = localMem[428];
              updateArrayLength(1, localMem[426], 5);
              ip = 955;
      end

        955 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 6] = 0;
              updateArrayLength(1, localMem[426], 6);
              ip = 956;
      end

        956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 3] = localMem[371];
              updateArrayLength(1, localMem[426], 3);
              ip = 957;
      end

        957 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[371]*6 + 1] = heapMem[localMem[371]*6 + 1] + 1;
              updateArrayLength(1, localMem[371], 1);
              ip = 958;
      end

        958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 1] = heapMem[localMem[371]*6 + 1];
              updateArrayLength(1, localMem[426], 1);
              ip = 959;
      end

        959 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[429] = !heapMem[localMem[360]*6 + 6];
              ip = 960;
      end

        960 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[429] != 0 ? 1012 : 961;
      end

        961 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[430] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[430] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[430]] = 0;
              ip = 962;
      end

        962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 6] = localMem[430];
              updateArrayLength(1, localMem[423], 6);
              ip = 963;
      end

        963 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[431] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[431] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[431]] = 0;
              ip = 964;
      end

        964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 6] = localMem[431];
              updateArrayLength(1, localMem[426], 6);
              ip = 965;
      end

        965 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[432] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 966;
      end

        966 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[433] = heapMem[localMem[423]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 967;
      end

        967 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[433] + 0 + i] = heapMem[NArea * localMem[432] + 0 + i];
                  updateArrayLength(1, localMem[433], 0 + i);
                end
              end
              ip = 968;
      end

        968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[434] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 969;
      end

        969 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[435] = heapMem[localMem[423]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 970;
      end

        970 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[435] + 0 + i] = heapMem[NArea * localMem[434] + 0 + i];
                  updateArrayLength(1, localMem[435], 0 + i);
                end
              end
              ip = 971;
      end

        971 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[436] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 972;
      end

        972 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[437] = heapMem[localMem[423]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 973;
      end

        973 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[438] = localMem[373] + 1;
              updateArrayLength(2, 0, 0);
              ip = 974;
      end

        974 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[438]) begin
                  heapMem[NArea * localMem[437] + 0 + i] = heapMem[NArea * localMem[436] + 0 + i];
                  updateArrayLength(1, localMem[437], 0 + i);
                end
              end
              ip = 975;
      end

        975 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[439] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 976;
      end

        976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[440] = heapMem[localMem[426]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 977;
      end

        977 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[440] + 0 + i] = heapMem[NArea * localMem[439] + localMem[374] + i];
                  updateArrayLength(1, localMem[440], 0 + i);
                end
              end
              ip = 978;
      end

        978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[441] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 979;
      end

        979 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[442] = heapMem[localMem[426]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 980;
      end

        980 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[442] + 0 + i] = heapMem[NArea * localMem[441] + localMem[374] + i];
                  updateArrayLength(1, localMem[442], 0 + i);
                end
              end
              ip = 981;
      end

        981 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[443] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 982;
      end

        982 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[444] = heapMem[localMem[426]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 983;
      end

        983 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[445] = localMem[373] + 1;
              updateArrayLength(2, 0, 0);
              ip = 984;
      end

        984 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[445]) begin
                  heapMem[NArea * localMem[444] + 0 + i] = heapMem[NArea * localMem[443] + localMem[374] + i];
                  updateArrayLength(1, localMem[444], 0 + i);
                end
              end
              ip = 985;
      end

        985 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[446] = heapMem[localMem[423]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 986;
      end

        986 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[447] = localMem[446] + 1;
              updateArrayLength(2, 0, 0);
              ip = 987;
      end

        987 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[448] = heapMem[localMem[423]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 988;
      end

        988 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 989;
      end

        989 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[449] = 0;
              updateArrayLength(2, 0, 0);
              ip = 990;
      end

        990 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 991;
      end

        991 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[449] >= localMem[447] ? 997 : 992;
      end

        992 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[450] = heapMem[localMem[448]*6 + localMem[449]];
              updateArrayLength(2, 0, 0);
              ip = 993;
      end

        993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[450]*6 + 2] = localMem[423];
              updateArrayLength(1, localMem[450], 2);
              ip = 994;
      end

        994 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 995;
      end

        995 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[449] = localMem[449] + 1;
              updateArrayLength(2, 0, 0);
              ip = 996;
      end

        996 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 990;
      end

        997 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 998;
      end

        998 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[451] = heapMem[localMem[426]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 999;
      end

        999 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[452] = localMem[451] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1000;
      end

       1000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[453] = heapMem[localMem[426]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1001;
      end

       1001 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1002;
      end

       1002 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[454] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1003;
      end

       1003 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1004;
      end

       1004 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[454] >= localMem[452] ? 1010 : 1005;
      end

       1005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[455] = heapMem[localMem[453]*6 + localMem[454]];
              updateArrayLength(2, 0, 0);
              ip = 1006;
      end

       1006 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[455]*6 + 2] = localMem[426];
              updateArrayLength(1, localMem[455], 2);
              ip = 1007;
      end

       1007 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1008;
      end

       1008 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[454] = localMem[454] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1009;
      end

       1009 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1003;
      end

       1010 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1011;
      end

       1011 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1027;
      end

       1012 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1013;
      end

       1013 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[456] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[456] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[456]] = 0;
              ip = 1014;
      end

       1014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[360]*6 + 6] = localMem[456];
              updateArrayLength(1, localMem[360], 6);
              ip = 1015;
      end

       1015 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[457] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1016;
      end

       1016 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[458] = heapMem[localMem[423]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1017;
      end

       1017 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[458] + 0 + i] = heapMem[NArea * localMem[457] + 0 + i];
                  updateArrayLength(1, localMem[458], 0 + i);
                end
              end
              ip = 1018;
      end

       1018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[459] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1019;
      end

       1019 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[460] = heapMem[localMem[423]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1020;
      end

       1020 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[460] + 0 + i] = heapMem[NArea * localMem[459] + 0 + i];
                  updateArrayLength(1, localMem[460], 0 + i);
                end
              end
              ip = 1021;
      end

       1021 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[461] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1022;
      end

       1022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[462] = heapMem[localMem[426]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1023;
      end

       1023 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[462] + 0 + i] = heapMem[NArea * localMem[461] + localMem[374] + i];
                  updateArrayLength(1, localMem[462], 0 + i);
                end
              end
              ip = 1024;
      end

       1024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[463] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1025;
      end

       1025 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[464] = heapMem[localMem[426]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1026;
      end

       1026 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[373]) begin
                  heapMem[NArea * localMem[464] + 0 + i] = heapMem[NArea * localMem[463] + localMem[374] + i];
                  updateArrayLength(1, localMem[464], 0 + i);
                end
              end
              ip = 1027;
      end

       1027 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1028;
      end

       1028 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[423]*6 + 2] = localMem[360];
              updateArrayLength(1, localMem[423], 2);
              ip = 1029;
      end

       1029 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[426]*6 + 2] = localMem[360];
              updateArrayLength(1, localMem[426], 2);
              ip = 1030;
      end

       1030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[465] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1031;
      end

       1031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[466] = heapMem[localMem[465]*6 + localMem[373]];
              updateArrayLength(2, 0, 0);
              ip = 1032;
      end

       1032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[467] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1033;
      end

       1033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[468] = heapMem[localMem[467]*6 + localMem[373]];
              updateArrayLength(2, 0, 0);
              ip = 1034;
      end

       1034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[469] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1035;
      end

       1035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[469]*6 + 0] = localMem[466];
              updateArrayLength(1, localMem[469], 0);
              ip = 1036;
      end

       1036 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[470] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1037;
      end

       1037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[470]*6 + 0] = localMem[468];
              updateArrayLength(1, localMem[470], 0);
              ip = 1038;
      end

       1038 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[471] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1039;
      end

       1039 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[471]*6 + 0] = localMem[423];
              updateArrayLength(1, localMem[471], 0);
              ip = 1040;
      end

       1040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[472] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1041;
      end

       1041 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[472]*6 + 1] = localMem[426];
              updateArrayLength(1, localMem[472], 1);
              ip = 1042;
      end

       1042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[360]*6 + 0] = 1;
              updateArrayLength(1, localMem[360], 0);
              ip = 1043;
      end

       1043 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[473] = heapMem[localMem[360]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1044;
      end

       1044 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[473]] = 1;
              ip = 1045;
      end

       1045 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[474] = heapMem[localMem[360]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1046;
      end

       1046 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[474]] = 1;
              ip = 1047;
      end

       1047 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[475] = heapMem[localMem[360]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1048;
      end

       1048 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[475]] = 2;
              ip = 1049;
      end

       1049 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1051;
      end

       1050 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1056;
      end

       1051 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1052;
      end

       1052 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[369] = 1;
              updateArrayLength(2, 0, 0);
              ip = 1053;
      end

       1053 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1056;
      end

       1054 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1055;
      end

       1055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[369] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1056;
      end

       1056 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1057;
      end

       1057 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1058;
      end

       1058 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1059;
      end

       1059 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1060;
      end

       1060 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[1]] = 0;
              freedArrays[freedArraysTop] = localMem[1];
              freedArraysTop = freedArraysTop + 1;
              ip = 1061;
      end

       1061 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[476] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[476] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[476]] = 0;
              ip = 1062;
      end

       1062 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1063;
      end

       1063 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[477] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1064;
      end

       1064 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[477] != 0 ? 1087 : 1065;
      end

       1065 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[478] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[478] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[478]] = 0;
              ip = 1066;
      end

       1066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 0] = 1;
              updateArrayLength(1, localMem[478], 0);
              ip = 1067;
      end

       1067 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 2] = 0;
              updateArrayLength(1, localMem[478], 2);
              ip = 1068;
      end

       1068 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[479] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[479] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[479]] = 0;
              ip = 1069;
      end

       1069 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 4] = localMem[479];
              updateArrayLength(1, localMem[478], 4);
              ip = 1070;
      end

       1070 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[480] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[480] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[480]] = 0;
              ip = 1071;
      end

       1071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 5] = localMem[480];
              updateArrayLength(1, localMem[478], 5);
              ip = 1072;
      end

       1072 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 6] = 0;
              updateArrayLength(1, localMem[478], 6);
              ip = 1073;
      end

       1073 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 3] = localMem[0];
              updateArrayLength(1, localMem[478], 3);
              ip = 1074;
      end

       1074 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = heapMem[localMem[0]*6 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 1075;
      end

       1075 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[478]*6 + 1] = heapMem[localMem[0]*6 + 1];
              updateArrayLength(1, localMem[478], 1);
              ip = 1076;
      end

       1076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[481] = heapMem[localMem[478]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1077;
      end

       1077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[481]*6 + 0] = 2;
              updateArrayLength(1, localMem[481], 0);
              ip = 1078;
      end

       1078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[482] = heapMem[localMem[478]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1079;
      end

       1079 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[482]*6 + 0] = 22;
              updateArrayLength(1, localMem[482], 0);
              ip = 1080;
      end

       1080 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 1081;
      end

       1081 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = localMem[478];
              updateArrayLength(1, localMem[0], 3);
              ip = 1082;
      end

       1082 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[483] = heapMem[localMem[478]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1083;
      end

       1083 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[483]] = 1;
              ip = 1084;
      end

       1084 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[484] = heapMem[localMem[478]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1085;
      end

       1085 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[484]] = 1;
              ip = 1086;
      end

       1086 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2115;
      end

       1087 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1088;
      end

       1088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[485] = heapMem[localMem[477]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1089;
      end

       1089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[486] = heapMem[localMem[0]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1090;
      end

       1090 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[485] >= localMem[486] ? 1126 : 1091;
      end

       1091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[487] = heapMem[localMem[477]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1092;
      end

       1092 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[487] != 0 ? 1125 : 1093;
      end

       1093 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[488] = !heapMem[localMem[477]*6 + 6];
              ip = 1094;
      end

       1094 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[488] == 0 ? 1124 : 1095;
      end

       1095 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[489] = heapMem[localMem[477]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1096;
      end

       1096 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[490] = 0; k = arraySizes[localMem[489]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[489] * NArea + i] == 2) localMem[490] = i + 1;
              end
              ip = 1097;
      end

       1097 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[490] == 0 ? 1102 : 1098;
      end

       1098 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[490] = localMem[490] - 1;
              updateArrayLength(2, 0, 0);
              ip = 1099;
      end

       1099 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[491] = heapMem[localMem[477]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1100;
      end

       1100 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[491]*6 + localMem[490]] = 22;
              updateArrayLength(1, localMem[491], localMem[490]);
              ip = 1101;
      end

       1101 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2115;
      end

       1102 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1103;
      end

       1103 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[489]] = localMem[485];
              ip = 1104;
      end

       1104 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[492] = heapMem[localMem[477]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1105;
      end

       1105 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[492]] = localMem[485];
              ip = 1106;
      end

       1106 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[489]];
//$display("AAAAA k=%d  source2=%d", k, 2);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[489] * NArea + i]);
                if (i < k && heapMem[localMem[489] * NArea + i] > 2) j = j + 1;
              end
              localMem[493] = j;
              ip = 1107;
      end

       1107 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[493] != 0 ? 1115 : 1108;
      end

       1108 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[494] = heapMem[localMem[477]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1109;
      end

       1109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[494]*6 + localMem[485]] = 2;
              updateArrayLength(1, localMem[494], localMem[485]);
              ip = 1110;
      end

       1110 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[495] = heapMem[localMem[477]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1111;
      end

       1111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[495]*6 + localMem[485]] = 22;
              updateArrayLength(1, localMem[495], localMem[485]);
              ip = 1112;
      end

       1112 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[477]*6 + 0] = localMem[485] + 1;
              updateArrayLength(1, localMem[477], 0);
              ip = 1113;
      end

       1113 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 1114;
      end

       1114 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2115;
      end

       1115 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1116;
      end

       1116 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[489]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[489] * NArea + i] < 2) j = j + 1;
              end
              localMem[496] = j;
              ip = 1117;
      end

       1117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[497] = heapMem[localMem[477]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1118;
      end

       1118 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[497] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[496], localMem[497], arraySizes[localMem[497]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[496] && i <= arraySizes[localMem[497]]) begin
                  heapMem[NArea * localMem[497] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[497] + localMem[496]] = 2;                                    // Insert new value
              arraySizes[localMem[497]] = arraySizes[localMem[497]] + 1;                              // Increase array size
              ip = 1119;
      end

       1119 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[498] = heapMem[localMem[477]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1120;
      end

       1120 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[498] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[496], localMem[498], arraySizes[localMem[498]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[496] && i <= arraySizes[localMem[498]]) begin
                  heapMem[NArea * localMem[498] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[498] + localMem[496]] = 22;                                    // Insert new value
              arraySizes[localMem[498]] = arraySizes[localMem[498]] + 1;                              // Increase array size
              ip = 1121;
      end

       1121 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[477]*6 + 0] = heapMem[localMem[477]*6 + 0] + 1;
              updateArrayLength(1, localMem[477], 0);
              ip = 1122;
      end

       1122 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 1123;
      end

       1123 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2115;
      end

       1124 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1125;
      end

       1125 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1126;
      end

       1126 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1127;
      end

       1127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[499] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1128;
      end

       1128 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1129;
      end

       1129 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[501] = heapMem[localMem[499]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1130;
      end

       1130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[502] = heapMem[localMem[499]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1131;
      end

       1131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[503] = heapMem[localMem[502]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1132;
      end

       1132 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[501] <  localMem[503] ? 1352 : 1133;
      end

       1133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[504] = localMem[503];
              updateArrayLength(2, 0, 0);
              ip = 1134;
      end

       1134 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[504] = localMem[504] >> 1;
              ip = 1135;
      end

       1135 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[505] = localMem[504] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1136;
      end

       1136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[506] = heapMem[localMem[499]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1137;
      end

       1137 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[506] == 0 ? 1234 : 1138;
      end

       1138 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[507] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[507] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[507]] = 0;
              ip = 1139;
      end

       1139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 0] = localMem[504];
              updateArrayLength(1, localMem[507], 0);
              ip = 1140;
      end

       1140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 2] = 0;
              updateArrayLength(1, localMem[507], 2);
              ip = 1141;
      end

       1141 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[508] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[508] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[508]] = 0;
              ip = 1142;
      end

       1142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 4] = localMem[508];
              updateArrayLength(1, localMem[507], 4);
              ip = 1143;
      end

       1143 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[509] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[509] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[509]] = 0;
              ip = 1144;
      end

       1144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 5] = localMem[509];
              updateArrayLength(1, localMem[507], 5);
              ip = 1145;
      end

       1145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 6] = 0;
              updateArrayLength(1, localMem[507], 6);
              ip = 1146;
      end

       1146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 3] = localMem[502];
              updateArrayLength(1, localMem[507], 3);
              ip = 1147;
      end

       1147 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[502]*6 + 1] = heapMem[localMem[502]*6 + 1] + 1;
              updateArrayLength(1, localMem[502], 1);
              ip = 1148;
      end

       1148 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 1] = heapMem[localMem[502]*6 + 1];
              updateArrayLength(1, localMem[507], 1);
              ip = 1149;
      end

       1149 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[510] = !heapMem[localMem[499]*6 + 6];
              ip = 1150;
      end

       1150 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[510] != 0 ? 1179 : 1151;
      end

       1151 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[511] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[511] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[511]] = 0;
              ip = 1152;
      end

       1152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 6] = localMem[511];
              updateArrayLength(1, localMem[507], 6);
              ip = 1153;
      end

       1153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[512] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1154;
      end

       1154 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[513] = heapMem[localMem[507]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1155;
      end

       1155 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[513] + 0 + i] = heapMem[NArea * localMem[512] + localMem[505] + i];
                  updateArrayLength(1, localMem[513], 0 + i);
                end
              end
              ip = 1156;
      end

       1156 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[514] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1157;
      end

       1157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[515] = heapMem[localMem[507]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1158;
      end

       1158 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[515] + 0 + i] = heapMem[NArea * localMem[514] + localMem[505] + i];
                  updateArrayLength(1, localMem[515], 0 + i);
                end
              end
              ip = 1159;
      end

       1159 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[516] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1160;
      end

       1160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[517] = heapMem[localMem[507]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1161;
      end

       1161 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[518] = localMem[504] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1162;
      end

       1162 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[518]) begin
                  heapMem[NArea * localMem[517] + 0 + i] = heapMem[NArea * localMem[516] + localMem[505] + i];
                  updateArrayLength(1, localMem[517], 0 + i);
                end
              end
              ip = 1163;
      end

       1163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[519] = heapMem[localMem[507]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1164;
      end

       1164 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[520] = localMem[519] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1165;
      end

       1165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[521] = heapMem[localMem[507]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1166;
      end

       1166 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1167;
      end

       1167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[522] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1168;
      end

       1168 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1169;
      end

       1169 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[522] >= localMem[520] ? 1175 : 1170;
      end

       1170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[523] = heapMem[localMem[521]*6 + localMem[522]];
              updateArrayLength(2, 0, 0);
              ip = 1171;
      end

       1171 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[523]*6 + 2] = localMem[507];
              updateArrayLength(1, localMem[523], 2);
              ip = 1172;
      end

       1172 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1173;
      end

       1173 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[522] = localMem[522] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1174;
      end

       1174 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1168;
      end

       1175 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1176;
      end

       1176 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[524] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1177;
      end

       1177 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[524]] = localMem[505];
              ip = 1178;
      end

       1178 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1186;
      end

       1179 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1180;
      end

       1180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[525] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1181;
      end

       1181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[526] = heapMem[localMem[507]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1182;
      end

       1182 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[526] + 0 + i] = heapMem[NArea * localMem[525] + localMem[505] + i];
                  updateArrayLength(1, localMem[526], 0 + i);
                end
              end
              ip = 1183;
      end

       1183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[527] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1184;
      end

       1184 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[528] = heapMem[localMem[507]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1185;
      end

       1185 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[528] + 0 + i] = heapMem[NArea * localMem[527] + localMem[505] + i];
                  updateArrayLength(1, localMem[528], 0 + i);
                end
              end
              ip = 1186;
      end

       1186 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1187;
      end

       1187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[499]*6 + 0] = localMem[504];
              updateArrayLength(1, localMem[499], 0);
              ip = 1188;
      end

       1188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[507]*6 + 2] = localMem[506];
              updateArrayLength(1, localMem[507], 2);
              ip = 1189;
      end

       1189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[529] = heapMem[localMem[506]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1190;
      end

       1190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[530] = heapMem[localMem[506]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1191;
      end

       1191 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[531] = heapMem[localMem[530]*6 + localMem[529]];
              updateArrayLength(2, 0, 0);
              ip = 1192;
      end

       1192 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[531] != localMem[499] ? 1211 : 1193;
      end

       1193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[532] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1194;
      end

       1194 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[533] = heapMem[localMem[532]*6 + localMem[504]];
              updateArrayLength(2, 0, 0);
              ip = 1195;
      end

       1195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[534] = heapMem[localMem[506]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1196;
      end

       1196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[534]*6 + localMem[529]] = localMem[533];
              updateArrayLength(1, localMem[534], localMem[529]);
              ip = 1197;
      end

       1197 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[535] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1198;
      end

       1198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[536] = heapMem[localMem[535]*6 + localMem[504]];
              updateArrayLength(2, 0, 0);
              ip = 1199;
      end

       1199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[537] = heapMem[localMem[506]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1200;
      end

       1200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[537]*6 + localMem[529]] = localMem[536];
              updateArrayLength(1, localMem[537], localMem[529]);
              ip = 1201;
      end

       1201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[538] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1202;
      end

       1202 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[538]] = localMem[504];
              ip = 1203;
      end

       1203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[539] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1204;
      end

       1204 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[539]] = localMem[504];
              ip = 1205;
      end

       1205 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[540] = localMem[529] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1206;
      end

       1206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[506]*6 + 0] = localMem[540];
              updateArrayLength(1, localMem[506], 0);
              ip = 1207;
      end

       1207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[541] = heapMem[localMem[506]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1208;
      end

       1208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[541]*6 + localMem[540]] = localMem[507];
              updateArrayLength(1, localMem[541], localMem[540]);
              ip = 1209;
      end

       1209 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1349;
      end

       1210 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1233;
      end

       1211 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1212;
      end

       1212 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 1213;
      end

       1213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[542] = heapMem[localMem[506]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1214;
      end

       1214 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[543] = 0; k = arraySizes[localMem[542]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[542] * NArea + i] == localMem[499]) localMem[543] = i + 1;
              end
              ip = 1215;
      end

       1215 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[543] = localMem[543] - 1;
              updateArrayLength(2, 0, 0);
              ip = 1216;
      end

       1216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[544] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1217;
      end

       1217 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[545] = heapMem[localMem[544]*6 + localMem[504]];
              updateArrayLength(2, 0, 0);
              ip = 1218;
      end

       1218 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[546] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1219;
      end

       1219 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[547] = heapMem[localMem[546]*6 + localMem[504]];
              updateArrayLength(2, 0, 0);
              ip = 1220;
      end

       1220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[548] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1221;
      end

       1221 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[548]] = localMem[504];
              ip = 1222;
      end

       1222 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[549] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1223;
      end

       1223 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[549]] = localMem[504];
              ip = 1224;
      end

       1224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[550] = heapMem[localMem[506]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1225;
      end

       1225 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[550] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[543], localMem[550], arraySizes[localMem[550]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[543] && i <= arraySizes[localMem[550]]) begin
                  heapMem[NArea * localMem[550] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[550] + localMem[543]] = localMem[545];                                    // Insert new value
              arraySizes[localMem[550]] = arraySizes[localMem[550]] + 1;                              // Increase array size
              ip = 1226;
      end

       1226 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[551] = heapMem[localMem[506]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1227;
      end

       1227 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[551] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[543], localMem[551], arraySizes[localMem[551]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[543] && i <= arraySizes[localMem[551]]) begin
                  heapMem[NArea * localMem[551] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[551] + localMem[543]] = localMem[547];                                    // Insert new value
              arraySizes[localMem[551]] = arraySizes[localMem[551]] + 1;                              // Increase array size
              ip = 1228;
      end

       1228 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[552] = heapMem[localMem[506]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1229;
      end

       1229 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[553] = localMem[543] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1230;
      end

       1230 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[552] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[553], localMem[552], arraySizes[localMem[552]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[553] && i <= arraySizes[localMem[552]]) begin
                  heapMem[NArea * localMem[552] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[552] + localMem[553]] = localMem[507];                                    // Insert new value
              arraySizes[localMem[552]] = arraySizes[localMem[552]] + 1;                              // Increase array size
              ip = 1231;
      end

       1231 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[506]*6 + 0] = heapMem[localMem[506]*6 + 0] + 1;
              updateArrayLength(1, localMem[506], 0);
              ip = 1232;
      end

       1232 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1349;
      end

       1233 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1234;
      end

       1234 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1235;
      end

       1235 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[554] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[554] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[554]] = 0;
              ip = 1236;
      end

       1236 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 0] = localMem[504];
              updateArrayLength(1, localMem[554], 0);
              ip = 1237;
      end

       1237 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 2] = 0;
              updateArrayLength(1, localMem[554], 2);
              ip = 1238;
      end

       1238 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[555] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[555] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[555]] = 0;
              ip = 1239;
      end

       1239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 4] = localMem[555];
              updateArrayLength(1, localMem[554], 4);
              ip = 1240;
      end

       1240 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[556] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[556] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[556]] = 0;
              ip = 1241;
      end

       1241 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 5] = localMem[556];
              updateArrayLength(1, localMem[554], 5);
              ip = 1242;
      end

       1242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 6] = 0;
              updateArrayLength(1, localMem[554], 6);
              ip = 1243;
      end

       1243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 3] = localMem[502];
              updateArrayLength(1, localMem[554], 3);
              ip = 1244;
      end

       1244 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[502]*6 + 1] = heapMem[localMem[502]*6 + 1] + 1;
              updateArrayLength(1, localMem[502], 1);
              ip = 1245;
      end

       1245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 1] = heapMem[localMem[502]*6 + 1];
              updateArrayLength(1, localMem[554], 1);
              ip = 1246;
      end

       1246 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[557] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[557] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[557]] = 0;
              ip = 1247;
      end

       1247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 0] = localMem[504];
              updateArrayLength(1, localMem[557], 0);
              ip = 1248;
      end

       1248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 2] = 0;
              updateArrayLength(1, localMem[557], 2);
              ip = 1249;
      end

       1249 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[558] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[558] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[558]] = 0;
              ip = 1250;
      end

       1250 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 4] = localMem[558];
              updateArrayLength(1, localMem[557], 4);
              ip = 1251;
      end

       1251 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[559] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[559] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[559]] = 0;
              ip = 1252;
      end

       1252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 5] = localMem[559];
              updateArrayLength(1, localMem[557], 5);
              ip = 1253;
      end

       1253 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 6] = 0;
              updateArrayLength(1, localMem[557], 6);
              ip = 1254;
      end

       1254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 3] = localMem[502];
              updateArrayLength(1, localMem[557], 3);
              ip = 1255;
      end

       1255 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[502]*6 + 1] = heapMem[localMem[502]*6 + 1] + 1;
              updateArrayLength(1, localMem[502], 1);
              ip = 1256;
      end

       1256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 1] = heapMem[localMem[502]*6 + 1];
              updateArrayLength(1, localMem[557], 1);
              ip = 1257;
      end

       1257 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[560] = !heapMem[localMem[499]*6 + 6];
              ip = 1258;
      end

       1258 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[560] != 0 ? 1310 : 1259;
      end

       1259 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[561] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[561] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[561]] = 0;
              ip = 1260;
      end

       1260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 6] = localMem[561];
              updateArrayLength(1, localMem[554], 6);
              ip = 1261;
      end

       1261 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[562] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[562] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[562]] = 0;
              ip = 1262;
      end

       1262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 6] = localMem[562];
              updateArrayLength(1, localMem[557], 6);
              ip = 1263;
      end

       1263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[563] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1264;
      end

       1264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[564] = heapMem[localMem[554]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1265;
      end

       1265 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[564] + 0 + i] = heapMem[NArea * localMem[563] + 0 + i];
                  updateArrayLength(1, localMem[564], 0 + i);
                end
              end
              ip = 1266;
      end

       1266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[565] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1267;
      end

       1267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[566] = heapMem[localMem[554]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1268;
      end

       1268 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[566] + 0 + i] = heapMem[NArea * localMem[565] + 0 + i];
                  updateArrayLength(1, localMem[566], 0 + i);
                end
              end
              ip = 1269;
      end

       1269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[567] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1270;
      end

       1270 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[568] = heapMem[localMem[554]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1271;
      end

       1271 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[569] = localMem[504] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1272;
      end

       1272 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[569]) begin
                  heapMem[NArea * localMem[568] + 0 + i] = heapMem[NArea * localMem[567] + 0 + i];
                  updateArrayLength(1, localMem[568], 0 + i);
                end
              end
              ip = 1273;
      end

       1273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[570] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1274;
      end

       1274 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[571] = heapMem[localMem[557]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1275;
      end

       1275 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[571] + 0 + i] = heapMem[NArea * localMem[570] + localMem[505] + i];
                  updateArrayLength(1, localMem[571], 0 + i);
                end
              end
              ip = 1276;
      end

       1276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[572] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1277;
      end

       1277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[573] = heapMem[localMem[557]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1278;
      end

       1278 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[573] + 0 + i] = heapMem[NArea * localMem[572] + localMem[505] + i];
                  updateArrayLength(1, localMem[573], 0 + i);
                end
              end
              ip = 1279;
      end

       1279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[574] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1280;
      end

       1280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[575] = heapMem[localMem[557]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1281;
      end

       1281 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[576] = localMem[504] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1282;
      end

       1282 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[576]) begin
                  heapMem[NArea * localMem[575] + 0 + i] = heapMem[NArea * localMem[574] + localMem[505] + i];
                  updateArrayLength(1, localMem[575], 0 + i);
                end
              end
              ip = 1283;
      end

       1283 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[577] = heapMem[localMem[554]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1284;
      end

       1284 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[578] = localMem[577] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1285;
      end

       1285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[579] = heapMem[localMem[554]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1286;
      end

       1286 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1287;
      end

       1287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[580] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1288;
      end

       1288 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1289;
      end

       1289 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[580] >= localMem[578] ? 1295 : 1290;
      end

       1290 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[581] = heapMem[localMem[579]*6 + localMem[580]];
              updateArrayLength(2, 0, 0);
              ip = 1291;
      end

       1291 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[581]*6 + 2] = localMem[554];
              updateArrayLength(1, localMem[581], 2);
              ip = 1292;
      end

       1292 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1293;
      end

       1293 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[580] = localMem[580] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1294;
      end

       1294 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1288;
      end

       1295 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1296;
      end

       1296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[582] = heapMem[localMem[557]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1297;
      end

       1297 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[583] = localMem[582] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1298;
      end

       1298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[584] = heapMem[localMem[557]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1299;
      end

       1299 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1300;
      end

       1300 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[585] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1301;
      end

       1301 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1302;
      end

       1302 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[585] >= localMem[583] ? 1308 : 1303;
      end

       1303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[586] = heapMem[localMem[584]*6 + localMem[585]];
              updateArrayLength(2, 0, 0);
              ip = 1304;
      end

       1304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[586]*6 + 2] = localMem[557];
              updateArrayLength(1, localMem[586], 2);
              ip = 1305;
      end

       1305 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1306;
      end

       1306 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[585] = localMem[585] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1307;
      end

       1307 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1301;
      end

       1308 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1309;
      end

       1309 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1325;
      end

       1310 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1311;
      end

       1311 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[587] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[587] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[587]] = 0;
              ip = 1312;
      end

       1312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[499]*6 + 6] = localMem[587];
              updateArrayLength(1, localMem[499], 6);
              ip = 1313;
      end

       1313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[588] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1314;
      end

       1314 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[589] = heapMem[localMem[554]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1315;
      end

       1315 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[589] + 0 + i] = heapMem[NArea * localMem[588] + 0 + i];
                  updateArrayLength(1, localMem[589], 0 + i);
                end
              end
              ip = 1316;
      end

       1316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[590] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1317;
      end

       1317 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[591] = heapMem[localMem[554]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1318;
      end

       1318 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[591] + 0 + i] = heapMem[NArea * localMem[590] + 0 + i];
                  updateArrayLength(1, localMem[591], 0 + i);
                end
              end
              ip = 1319;
      end

       1319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[592] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1320;
      end

       1320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[593] = heapMem[localMem[557]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1321;
      end

       1321 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[593] + 0 + i] = heapMem[NArea * localMem[592] + localMem[505] + i];
                  updateArrayLength(1, localMem[593], 0 + i);
                end
              end
              ip = 1322;
      end

       1322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[594] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1323;
      end

       1323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[595] = heapMem[localMem[557]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1324;
      end

       1324 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[504]) begin
                  heapMem[NArea * localMem[595] + 0 + i] = heapMem[NArea * localMem[594] + localMem[505] + i];
                  updateArrayLength(1, localMem[595], 0 + i);
                end
              end
              ip = 1325;
      end

       1325 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1326;
      end

       1326 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[554]*6 + 2] = localMem[499];
              updateArrayLength(1, localMem[554], 2);
              ip = 1327;
      end

       1327 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[557]*6 + 2] = localMem[499];
              updateArrayLength(1, localMem[557], 2);
              ip = 1328;
      end

       1328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[596] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1329;
      end

       1329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[597] = heapMem[localMem[596]*6 + localMem[504]];
              updateArrayLength(2, 0, 0);
              ip = 1330;
      end

       1330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[598] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1331;
      end

       1331 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[599] = heapMem[localMem[598]*6 + localMem[504]];
              updateArrayLength(2, 0, 0);
              ip = 1332;
      end

       1332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[600] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1333;
      end

       1333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[600]*6 + 0] = localMem[597];
              updateArrayLength(1, localMem[600], 0);
              ip = 1334;
      end

       1334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[601] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1335;
      end

       1335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[601]*6 + 0] = localMem[599];
              updateArrayLength(1, localMem[601], 0);
              ip = 1336;
      end

       1336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[602] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1337;
      end

       1337 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[602]*6 + 0] = localMem[554];
              updateArrayLength(1, localMem[602], 0);
              ip = 1338;
      end

       1338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[603] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1339;
      end

       1339 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[603]*6 + 1] = localMem[557];
              updateArrayLength(1, localMem[603], 1);
              ip = 1340;
      end

       1340 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[499]*6 + 0] = 1;
              updateArrayLength(1, localMem[499], 0);
              ip = 1341;
      end

       1341 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[604] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1342;
      end

       1342 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[604]] = 1;
              ip = 1343;
      end

       1343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[605] = heapMem[localMem[499]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1344;
      end

       1344 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[605]] = 1;
              ip = 1345;
      end

       1345 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[606] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1346;
      end

       1346 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[606]] = 2;
              ip = 1347;
      end

       1347 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1349;
      end

       1348 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1354;
      end

       1349 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1350;
      end

       1350 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[500] = 1;
              updateArrayLength(2, 0, 0);
              ip = 1351;
      end

       1351 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1354;
      end

       1352 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1353;
      end

       1353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[500] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1354;
      end

       1354 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1355;
      end

       1355 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1356;
      end

       1356 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1357;
      end

       1357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[607] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1358;
      end

       1358 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1359;
      end

       1359 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[607] >= 99 ? 1857 : 1360;
      end

       1360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[608] = heapMem[localMem[499]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1361;
      end

       1361 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[609] = localMem[608] - 1;
              updateArrayLength(2, 0, 0);
              ip = 1362;
      end

       1362 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[610] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1363;
      end

       1363 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[611] = heapMem[localMem[610]*6 + localMem[609]];
              updateArrayLength(2, 0, 0);
              ip = 1364;
      end

       1364 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 2 <= localMem[611] ? 1605 : 1365;
      end

       1365 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[612] = !heapMem[localMem[499]*6 + 6];
              ip = 1366;
      end

       1366 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[612] == 0 ? 1371 : 1367;
      end

       1367 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 0] = localMem[499];
              updateArrayLength(1, localMem[476], 0);
              ip = 1368;
      end

       1368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 1] = 2;
              updateArrayLength(1, localMem[476], 1);
              ip = 1369;
      end

       1369 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[476]*6 + 2] = localMem[608] - 1;
              updateArrayLength(1, localMem[476], 2);
              ip = 1370;
      end

       1370 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1861;
      end

       1371 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1372;
      end

       1372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[613] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1373;
      end

       1373 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[614] = heapMem[localMem[613]*6 + localMem[608]];
              updateArrayLength(2, 0, 0);
              ip = 1374;
      end

       1374 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1375;
      end

       1375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[616] = heapMem[localMem[614]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1376;
      end

       1376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[617] = heapMem[localMem[614]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1377;
      end

       1377 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[618] = heapMem[localMem[617]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1378;
      end

       1378 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[616] <  localMem[618] ? 1598 : 1379;
      end

       1379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[619] = localMem[618];
              updateArrayLength(2, 0, 0);
              ip = 1380;
      end

       1380 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[619] = localMem[619] >> 1;
              ip = 1381;
      end

       1381 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[620] = localMem[619] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1382;
      end

       1382 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[621] = heapMem[localMem[614]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1383;
      end

       1383 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[621] == 0 ? 1480 : 1384;
      end

       1384 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[622] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[622] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[622]] = 0;
              ip = 1385;
      end

       1385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 0] = localMem[619];
              updateArrayLength(1, localMem[622], 0);
              ip = 1386;
      end

       1386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 2] = 0;
              updateArrayLength(1, localMem[622], 2);
              ip = 1387;
      end

       1387 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[623] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[623] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[623]] = 0;
              ip = 1388;
      end

       1388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 4] = localMem[623];
              updateArrayLength(1, localMem[622], 4);
              ip = 1389;
      end

       1389 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[624] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[624] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[624]] = 0;
              ip = 1390;
      end

       1390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 5] = localMem[624];
              updateArrayLength(1, localMem[622], 5);
              ip = 1391;
      end

       1391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 6] = 0;
              updateArrayLength(1, localMem[622], 6);
              ip = 1392;
      end

       1392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 3] = localMem[617];
              updateArrayLength(1, localMem[622], 3);
              ip = 1393;
      end

       1393 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[617]*6 + 1] = heapMem[localMem[617]*6 + 1] + 1;
              updateArrayLength(1, localMem[617], 1);
              ip = 1394;
      end

       1394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 1] = heapMem[localMem[617]*6 + 1];
              updateArrayLength(1, localMem[622], 1);
              ip = 1395;
      end

       1395 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[625] = !heapMem[localMem[614]*6 + 6];
              ip = 1396;
      end

       1396 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[625] != 0 ? 1425 : 1397;
      end

       1397 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[626] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[626] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[626]] = 0;
              ip = 1398;
      end

       1398 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 6] = localMem[626];
              updateArrayLength(1, localMem[622], 6);
              ip = 1399;
      end

       1399 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[627] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1400;
      end

       1400 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[628] = heapMem[localMem[622]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1401;
      end

       1401 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[628] + 0 + i] = heapMem[NArea * localMem[627] + localMem[620] + i];
                  updateArrayLength(1, localMem[628], 0 + i);
                end
              end
              ip = 1402;
      end

       1402 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[629] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1403;
      end

       1403 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[630] = heapMem[localMem[622]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1404;
      end

       1404 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[630] + 0 + i] = heapMem[NArea * localMem[629] + localMem[620] + i];
                  updateArrayLength(1, localMem[630], 0 + i);
                end
              end
              ip = 1405;
      end

       1405 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[631] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1406;
      end

       1406 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[632] = heapMem[localMem[622]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1407;
      end

       1407 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[633] = localMem[619] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1408;
      end

       1408 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[633]) begin
                  heapMem[NArea * localMem[632] + 0 + i] = heapMem[NArea * localMem[631] + localMem[620] + i];
                  updateArrayLength(1, localMem[632], 0 + i);
                end
              end
              ip = 1409;
      end

       1409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[634] = heapMem[localMem[622]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1410;
      end

       1410 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[635] = localMem[634] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1411;
      end

       1411 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[636] = heapMem[localMem[622]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1412;
      end

       1412 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1413;
      end

       1413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[637] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1414;
      end

       1414 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1415;
      end

       1415 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[637] >= localMem[635] ? 1421 : 1416;
      end

       1416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[638] = heapMem[localMem[636]*6 + localMem[637]];
              updateArrayLength(2, 0, 0);
              ip = 1417;
      end

       1417 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[638]*6 + 2] = localMem[622];
              updateArrayLength(1, localMem[638], 2);
              ip = 1418;
      end

       1418 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1419;
      end

       1419 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[637] = localMem[637] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1420;
      end

       1420 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1414;
      end

       1421 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1422;
      end

       1422 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[639] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1423;
      end

       1423 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[639]] = localMem[620];
              ip = 1424;
      end

       1424 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1432;
      end

       1425 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1426;
      end

       1426 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[640] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1427;
      end

       1427 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[641] = heapMem[localMem[622]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1428;
      end

       1428 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[641] + 0 + i] = heapMem[NArea * localMem[640] + localMem[620] + i];
                  updateArrayLength(1, localMem[641], 0 + i);
                end
              end
              ip = 1429;
      end

       1429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[642] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1430;
      end

       1430 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[643] = heapMem[localMem[622]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1431;
      end

       1431 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[643] + 0 + i] = heapMem[NArea * localMem[642] + localMem[620] + i];
                  updateArrayLength(1, localMem[643], 0 + i);
                end
              end
              ip = 1432;
      end

       1432 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1433;
      end

       1433 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[614]*6 + 0] = localMem[619];
              updateArrayLength(1, localMem[614], 0);
              ip = 1434;
      end

       1434 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[622]*6 + 2] = localMem[621];
              updateArrayLength(1, localMem[622], 2);
              ip = 1435;
      end

       1435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[644] = heapMem[localMem[621]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1436;
      end

       1436 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[645] = heapMem[localMem[621]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1437;
      end

       1437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[646] = heapMem[localMem[645]*6 + localMem[644]];
              updateArrayLength(2, 0, 0);
              ip = 1438;
      end

       1438 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[646] != localMem[614] ? 1457 : 1439;
      end

       1439 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[647] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1440;
      end

       1440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[648] = heapMem[localMem[647]*6 + localMem[619]];
              updateArrayLength(2, 0, 0);
              ip = 1441;
      end

       1441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[649] = heapMem[localMem[621]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1442;
      end

       1442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[649]*6 + localMem[644]] = localMem[648];
              updateArrayLength(1, localMem[649], localMem[644]);
              ip = 1443;
      end

       1443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[650] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1444;
      end

       1444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[651] = heapMem[localMem[650]*6 + localMem[619]];
              updateArrayLength(2, 0, 0);
              ip = 1445;
      end

       1445 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[652] = heapMem[localMem[621]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1446;
      end

       1446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[652]*6 + localMem[644]] = localMem[651];
              updateArrayLength(1, localMem[652], localMem[644]);
              ip = 1447;
      end

       1447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[653] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1448;
      end

       1448 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[653]] = localMem[619];
              ip = 1449;
      end

       1449 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[654] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1450;
      end

       1450 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[654]] = localMem[619];
              ip = 1451;
      end

       1451 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[655] = localMem[644] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1452;
      end

       1452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[621]*6 + 0] = localMem[655];
              updateArrayLength(1, localMem[621], 0);
              ip = 1453;
      end

       1453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[656] = heapMem[localMem[621]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1454;
      end

       1454 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[656]*6 + localMem[655]] = localMem[622];
              updateArrayLength(1, localMem[656], localMem[655]);
              ip = 1455;
      end

       1455 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1595;
      end

       1456 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1479;
      end

       1457 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1458;
      end

       1458 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 1459;
      end

       1459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[657] = heapMem[localMem[621]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1460;
      end

       1460 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[658] = 0; k = arraySizes[localMem[657]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[657] * NArea + i] == localMem[614]) localMem[658] = i + 1;
              end
              ip = 1461;
      end

       1461 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[658] = localMem[658] - 1;
              updateArrayLength(2, 0, 0);
              ip = 1462;
      end

       1462 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[659] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1463;
      end

       1463 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[660] = heapMem[localMem[659]*6 + localMem[619]];
              updateArrayLength(2, 0, 0);
              ip = 1464;
      end

       1464 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[661] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1465;
      end

       1465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[662] = heapMem[localMem[661]*6 + localMem[619]];
              updateArrayLength(2, 0, 0);
              ip = 1466;
      end

       1466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[663] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1467;
      end

       1467 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[663]] = localMem[619];
              ip = 1468;
      end

       1468 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[664] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1469;
      end

       1469 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[664]] = localMem[619];
              ip = 1470;
      end

       1470 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[665] = heapMem[localMem[621]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1471;
      end

       1471 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[665] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[658], localMem[665], arraySizes[localMem[665]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[658] && i <= arraySizes[localMem[665]]) begin
                  heapMem[NArea * localMem[665] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[665] + localMem[658]] = localMem[660];                                    // Insert new value
              arraySizes[localMem[665]] = arraySizes[localMem[665]] + 1;                              // Increase array size
              ip = 1472;
      end

       1472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[666] = heapMem[localMem[621]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1473;
      end

       1473 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[666] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[658], localMem[666], arraySizes[localMem[666]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[658] && i <= arraySizes[localMem[666]]) begin
                  heapMem[NArea * localMem[666] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[666] + localMem[658]] = localMem[662];                                    // Insert new value
              arraySizes[localMem[666]] = arraySizes[localMem[666]] + 1;                              // Increase array size
              ip = 1474;
      end

       1474 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[667] = heapMem[localMem[621]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1475;
      end

       1475 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[668] = localMem[658] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1476;
      end

       1476 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[667] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[668], localMem[667], arraySizes[localMem[667]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[668] && i <= arraySizes[localMem[667]]) begin
                  heapMem[NArea * localMem[667] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[667] + localMem[668]] = localMem[622];                                    // Insert new value
              arraySizes[localMem[667]] = arraySizes[localMem[667]] + 1;                              // Increase array size
              ip = 1477;
      end

       1477 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[621]*6 + 0] = heapMem[localMem[621]*6 + 0] + 1;
              updateArrayLength(1, localMem[621], 0);
              ip = 1478;
      end

       1478 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1595;
      end

       1479 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1480;
      end

       1480 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1481;
      end

       1481 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[669] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[669] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[669]] = 0;
              ip = 1482;
      end

       1482 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 0] = localMem[619];
              updateArrayLength(1, localMem[669], 0);
              ip = 1483;
      end

       1483 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 2] = 0;
              updateArrayLength(1, localMem[669], 2);
              ip = 1484;
      end

       1484 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[670] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[670] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[670]] = 0;
              ip = 1485;
      end

       1485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 4] = localMem[670];
              updateArrayLength(1, localMem[669], 4);
              ip = 1486;
      end

       1486 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[671] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[671] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[671]] = 0;
              ip = 1487;
      end

       1487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 5] = localMem[671];
              updateArrayLength(1, localMem[669], 5);
              ip = 1488;
      end

       1488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 6] = 0;
              updateArrayLength(1, localMem[669], 6);
              ip = 1489;
      end

       1489 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 3] = localMem[617];
              updateArrayLength(1, localMem[669], 3);
              ip = 1490;
      end

       1490 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[617]*6 + 1] = heapMem[localMem[617]*6 + 1] + 1;
              updateArrayLength(1, localMem[617], 1);
              ip = 1491;
      end

       1491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 1] = heapMem[localMem[617]*6 + 1];
              updateArrayLength(1, localMem[669], 1);
              ip = 1492;
      end

       1492 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[672] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[672] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[672]] = 0;
              ip = 1493;
      end

       1493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 0] = localMem[619];
              updateArrayLength(1, localMem[672], 0);
              ip = 1494;
      end

       1494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 2] = 0;
              updateArrayLength(1, localMem[672], 2);
              ip = 1495;
      end

       1495 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[673] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[673] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[673]] = 0;
              ip = 1496;
      end

       1496 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 4] = localMem[673];
              updateArrayLength(1, localMem[672], 4);
              ip = 1497;
      end

       1497 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[674] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[674] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[674]] = 0;
              ip = 1498;
      end

       1498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 5] = localMem[674];
              updateArrayLength(1, localMem[672], 5);
              ip = 1499;
      end

       1499 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 6] = 0;
              updateArrayLength(1, localMem[672], 6);
              ip = 1500;
      end

       1500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 3] = localMem[617];
              updateArrayLength(1, localMem[672], 3);
              ip = 1501;
      end

       1501 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[617]*6 + 1] = heapMem[localMem[617]*6 + 1] + 1;
              updateArrayLength(1, localMem[617], 1);
              ip = 1502;
      end

       1502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 1] = heapMem[localMem[617]*6 + 1];
              updateArrayLength(1, localMem[672], 1);
              ip = 1503;
      end

       1503 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[675] = !heapMem[localMem[614]*6 + 6];
              ip = 1504;
      end

       1504 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[675] != 0 ? 1556 : 1505;
      end

       1505 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[676] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[676] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[676]] = 0;
              ip = 1506;
      end

       1506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 6] = localMem[676];
              updateArrayLength(1, localMem[669], 6);
              ip = 1507;
      end

       1507 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[677] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[677] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[677]] = 0;
              ip = 1508;
      end

       1508 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 6] = localMem[677];
              updateArrayLength(1, localMem[672], 6);
              ip = 1509;
      end

       1509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[678] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1510;
      end

       1510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[679] = heapMem[localMem[669]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1511;
      end

       1511 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[679] + 0 + i] = heapMem[NArea * localMem[678] + 0 + i];
                  updateArrayLength(1, localMem[679], 0 + i);
                end
              end
              ip = 1512;
      end

       1512 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[680] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1513;
      end

       1513 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[681] = heapMem[localMem[669]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1514;
      end

       1514 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[681] + 0 + i] = heapMem[NArea * localMem[680] + 0 + i];
                  updateArrayLength(1, localMem[681], 0 + i);
                end
              end
              ip = 1515;
      end

       1515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[682] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1516;
      end

       1516 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[683] = heapMem[localMem[669]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1517;
      end

       1517 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[684] = localMem[619] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1518;
      end

       1518 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[684]) begin
                  heapMem[NArea * localMem[683] + 0 + i] = heapMem[NArea * localMem[682] + 0 + i];
                  updateArrayLength(1, localMem[683], 0 + i);
                end
              end
              ip = 1519;
      end

       1519 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[685] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1520;
      end

       1520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[686] = heapMem[localMem[672]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1521;
      end

       1521 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[686] + 0 + i] = heapMem[NArea * localMem[685] + localMem[620] + i];
                  updateArrayLength(1, localMem[686], 0 + i);
                end
              end
              ip = 1522;
      end

       1522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[687] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1523;
      end

       1523 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[688] = heapMem[localMem[672]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1524;
      end

       1524 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[688] + 0 + i] = heapMem[NArea * localMem[687] + localMem[620] + i];
                  updateArrayLength(1, localMem[688], 0 + i);
                end
              end
              ip = 1525;
      end

       1525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[689] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1526;
      end

       1526 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[690] = heapMem[localMem[672]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1527;
      end

       1527 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[691] = localMem[619] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1528;
      end

       1528 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[691]) begin
                  heapMem[NArea * localMem[690] + 0 + i] = heapMem[NArea * localMem[689] + localMem[620] + i];
                  updateArrayLength(1, localMem[690], 0 + i);
                end
              end
              ip = 1529;
      end

       1529 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[692] = heapMem[localMem[669]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1530;
      end

       1530 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[693] = localMem[692] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1531;
      end

       1531 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[694] = heapMem[localMem[669]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1532;
      end

       1532 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1533;
      end

       1533 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[695] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1534;
      end

       1534 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1535;
      end

       1535 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[695] >= localMem[693] ? 1541 : 1536;
      end

       1536 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[696] = heapMem[localMem[694]*6 + localMem[695]];
              updateArrayLength(2, 0, 0);
              ip = 1537;
      end

       1537 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[696]*6 + 2] = localMem[669];
              updateArrayLength(1, localMem[696], 2);
              ip = 1538;
      end

       1538 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1539;
      end

       1539 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[695] = localMem[695] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1540;
      end

       1540 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1534;
      end

       1541 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1542;
      end

       1542 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[697] = heapMem[localMem[672]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1543;
      end

       1543 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[698] = localMem[697] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1544;
      end

       1544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[699] = heapMem[localMem[672]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1545;
      end

       1545 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1546;
      end

       1546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[700] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1547;
      end

       1547 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1548;
      end

       1548 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[700] >= localMem[698] ? 1554 : 1549;
      end

       1549 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[701] = heapMem[localMem[699]*6 + localMem[700]];
              updateArrayLength(2, 0, 0);
              ip = 1550;
      end

       1550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[701]*6 + 2] = localMem[672];
              updateArrayLength(1, localMem[701], 2);
              ip = 1551;
      end

       1551 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1552;
      end

       1552 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[700] = localMem[700] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1553;
      end

       1553 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1547;
      end

       1554 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1555;
      end

       1555 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1571;
      end

       1556 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1557;
      end

       1557 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[702] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[702] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[702]] = 0;
              ip = 1558;
      end

       1558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[614]*6 + 6] = localMem[702];
              updateArrayLength(1, localMem[614], 6);
              ip = 1559;
      end

       1559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[703] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1560;
      end

       1560 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[704] = heapMem[localMem[669]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1561;
      end

       1561 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[704] + 0 + i] = heapMem[NArea * localMem[703] + 0 + i];
                  updateArrayLength(1, localMem[704], 0 + i);
                end
              end
              ip = 1562;
      end

       1562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[705] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1563;
      end

       1563 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[706] = heapMem[localMem[669]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1564;
      end

       1564 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[706] + 0 + i] = heapMem[NArea * localMem[705] + 0 + i];
                  updateArrayLength(1, localMem[706], 0 + i);
                end
              end
              ip = 1565;
      end

       1565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[707] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1566;
      end

       1566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[708] = heapMem[localMem[672]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1567;
      end

       1567 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[708] + 0 + i] = heapMem[NArea * localMem[707] + localMem[620] + i];
                  updateArrayLength(1, localMem[708], 0 + i);
                end
              end
              ip = 1568;
      end

       1568 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[709] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1569;
      end

       1569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[710] = heapMem[localMem[672]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1570;
      end

       1570 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[619]) begin
                  heapMem[NArea * localMem[710] + 0 + i] = heapMem[NArea * localMem[709] + localMem[620] + i];
                  updateArrayLength(1, localMem[710], 0 + i);
                end
              end
              ip = 1571;
      end

       1571 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1572;
      end

       1572 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[669]*6 + 2] = localMem[614];
              updateArrayLength(1, localMem[669], 2);
              ip = 1573;
      end

       1573 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[672]*6 + 2] = localMem[614];
              updateArrayLength(1, localMem[672], 2);
              ip = 1574;
      end

       1574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[711] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1575;
      end

       1575 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[712] = heapMem[localMem[711]*6 + localMem[619]];
              updateArrayLength(2, 0, 0);
              ip = 1576;
      end

       1576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[713] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1577;
      end

       1577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[714] = heapMem[localMem[713]*6 + localMem[619]];
              updateArrayLength(2, 0, 0);
              ip = 1578;
      end

       1578 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[715] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1579;
      end

       1579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[715]*6 + 0] = localMem[712];
              updateArrayLength(1, localMem[715], 0);
              ip = 1580;
      end

       1580 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[716] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1581;
      end

       1581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[716]*6 + 0] = localMem[714];
              updateArrayLength(1, localMem[716], 0);
              ip = 1582;
      end

       1582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[717] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1583;
      end

       1583 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[717]*6 + 0] = localMem[669];
              updateArrayLength(1, localMem[717], 0);
              ip = 1584;
      end

       1584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[718] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1585;
      end

       1585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[718]*6 + 1] = localMem[672];
              updateArrayLength(1, localMem[718], 1);
              ip = 1586;
      end

       1586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[614]*6 + 0] = 1;
              updateArrayLength(1, localMem[614], 0);
              ip = 1587;
      end

       1587 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[719] = heapMem[localMem[614]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1588;
      end

       1588 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[719]] = 1;
              ip = 1589;
      end

       1589 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[720] = heapMem[localMem[614]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1590;
      end

       1590 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[720]] = 1;
              ip = 1591;
      end

       1591 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[721] = heapMem[localMem[614]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1592;
      end

       1592 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[721]] = 2;
              ip = 1593;
      end

       1593 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1595;
      end

       1594 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1600;
      end

       1595 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1596;
      end

       1596 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[615] = 1;
              updateArrayLength(2, 0, 0);
              ip = 1597;
      end

       1597 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1600;
      end

       1598 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1599;
      end

       1599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[615] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1600;
      end

       1600 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1601;
      end

       1601 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[615] != 0 ? 1603 : 1602;
      end

       1602 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[499] = localMem[614];
              updateArrayLength(2, 0, 0);
              ip = 1603;
      end

       1603 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1604;
      end

       1604 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1854;
      end

       1605 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1606;
      end

       1606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[722] = heapMem[localMem[499]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1607;
      end

       1607 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[723] = 0; k = arraySizes[localMem[722]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[722] * NArea + i] == 2) localMem[723] = i + 1;
              end
              ip = 1608;
      end

       1608 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[723] == 0 ? 1613 : 1609;
      end

       1609 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 0] = localMem[499];
              updateArrayLength(1, localMem[476], 0);
              ip = 1610;
      end

       1610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 1] = 1;
              updateArrayLength(1, localMem[476], 1);
              ip = 1611;
      end

       1611 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[476]*6 + 2] = localMem[723] - 1;
              updateArrayLength(1, localMem[476], 2);
              ip = 1612;
      end

       1612 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1861;
      end

       1613 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1614;
      end

       1614 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[722]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[722] * NArea + i] < 2) j = j + 1;
              end
              localMem[724] = j;
              ip = 1615;
      end

       1615 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[725] = !heapMem[localMem[499]*6 + 6];
              ip = 1616;
      end

       1616 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[725] == 0 ? 1621 : 1617;
      end

       1617 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 0] = localMem[499];
              updateArrayLength(1, localMem[476], 0);
              ip = 1618;
      end

       1618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 1] = 0;
              updateArrayLength(1, localMem[476], 1);
              ip = 1619;
      end

       1619 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[476]*6 + 2] = localMem[724];
              updateArrayLength(1, localMem[476], 2);
              ip = 1620;
      end

       1620 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1861;
      end

       1621 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1622;
      end

       1622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[726] = heapMem[localMem[499]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1623;
      end

       1623 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[727] = heapMem[localMem[726]*6 + localMem[724]];
              updateArrayLength(2, 0, 0);
              ip = 1624;
      end

       1624 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1625;
      end

       1625 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[729] = heapMem[localMem[727]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1626;
      end

       1626 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[730] = heapMem[localMem[727]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1627;
      end

       1627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[731] = heapMem[localMem[730]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1628;
      end

       1628 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[729] <  localMem[731] ? 1848 : 1629;
      end

       1629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[732] = localMem[731];
              updateArrayLength(2, 0, 0);
              ip = 1630;
      end

       1630 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[732] = localMem[732] >> 1;
              ip = 1631;
      end

       1631 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[733] = localMem[732] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1632;
      end

       1632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[734] = heapMem[localMem[727]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1633;
      end

       1633 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[734] == 0 ? 1730 : 1634;
      end

       1634 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[735] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[735] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[735]] = 0;
              ip = 1635;
      end

       1635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 0] = localMem[732];
              updateArrayLength(1, localMem[735], 0);
              ip = 1636;
      end

       1636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 2] = 0;
              updateArrayLength(1, localMem[735], 2);
              ip = 1637;
      end

       1637 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[736] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[736] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[736]] = 0;
              ip = 1638;
      end

       1638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 4] = localMem[736];
              updateArrayLength(1, localMem[735], 4);
              ip = 1639;
      end

       1639 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[737] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[737] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[737]] = 0;
              ip = 1640;
      end

       1640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 5] = localMem[737];
              updateArrayLength(1, localMem[735], 5);
              ip = 1641;
      end

       1641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 6] = 0;
              updateArrayLength(1, localMem[735], 6);
              ip = 1642;
      end

       1642 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 3] = localMem[730];
              updateArrayLength(1, localMem[735], 3);
              ip = 1643;
      end

       1643 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[730]*6 + 1] = heapMem[localMem[730]*6 + 1] + 1;
              updateArrayLength(1, localMem[730], 1);
              ip = 1644;
      end

       1644 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 1] = heapMem[localMem[730]*6 + 1];
              updateArrayLength(1, localMem[735], 1);
              ip = 1645;
      end

       1645 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[738] = !heapMem[localMem[727]*6 + 6];
              ip = 1646;
      end

       1646 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[738] != 0 ? 1675 : 1647;
      end

       1647 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[739] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[739] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[739]] = 0;
              ip = 1648;
      end

       1648 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 6] = localMem[739];
              updateArrayLength(1, localMem[735], 6);
              ip = 1649;
      end

       1649 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[740] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1650;
      end

       1650 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[741] = heapMem[localMem[735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1651;
      end

       1651 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[741] + 0 + i] = heapMem[NArea * localMem[740] + localMem[733] + i];
                  updateArrayLength(1, localMem[741], 0 + i);
                end
              end
              ip = 1652;
      end

       1652 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[742] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1653;
      end

       1653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[743] = heapMem[localMem[735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1654;
      end

       1654 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[743] + 0 + i] = heapMem[NArea * localMem[742] + localMem[733] + i];
                  updateArrayLength(1, localMem[743], 0 + i);
                end
              end
              ip = 1655;
      end

       1655 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[744] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1656;
      end

       1656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[745] = heapMem[localMem[735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1657;
      end

       1657 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[746] = localMem[732] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1658;
      end

       1658 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[746]) begin
                  heapMem[NArea * localMem[745] + 0 + i] = heapMem[NArea * localMem[744] + localMem[733] + i];
                  updateArrayLength(1, localMem[745], 0 + i);
                end
              end
              ip = 1659;
      end

       1659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[747] = heapMem[localMem[735]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1660;
      end

       1660 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[748] = localMem[747] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1661;
      end

       1661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[749] = heapMem[localMem[735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1662;
      end

       1662 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1663;
      end

       1663 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[750] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1664;
      end

       1664 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1665;
      end

       1665 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[750] >= localMem[748] ? 1671 : 1666;
      end

       1666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[751] = heapMem[localMem[749]*6 + localMem[750]];
              updateArrayLength(2, 0, 0);
              ip = 1667;
      end

       1667 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[751]*6 + 2] = localMem[735];
              updateArrayLength(1, localMem[751], 2);
              ip = 1668;
      end

       1668 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1669;
      end

       1669 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[750] = localMem[750] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1670;
      end

       1670 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1664;
      end

       1671 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1672;
      end

       1672 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[752] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1673;
      end

       1673 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[752]] = localMem[733];
              ip = 1674;
      end

       1674 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1682;
      end

       1675 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1676;
      end

       1676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[753] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1677;
      end

       1677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[754] = heapMem[localMem[735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1678;
      end

       1678 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[754] + 0 + i] = heapMem[NArea * localMem[753] + localMem[733] + i];
                  updateArrayLength(1, localMem[754], 0 + i);
                end
              end
              ip = 1679;
      end

       1679 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[755] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1680;
      end

       1680 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[756] = heapMem[localMem[735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1681;
      end

       1681 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[756] + 0 + i] = heapMem[NArea * localMem[755] + localMem[733] + i];
                  updateArrayLength(1, localMem[756], 0 + i);
                end
              end
              ip = 1682;
      end

       1682 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1683;
      end

       1683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[727]*6 + 0] = localMem[732];
              updateArrayLength(1, localMem[727], 0);
              ip = 1684;
      end

       1684 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[735]*6 + 2] = localMem[734];
              updateArrayLength(1, localMem[735], 2);
              ip = 1685;
      end

       1685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[757] = heapMem[localMem[734]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1686;
      end

       1686 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[758] = heapMem[localMem[734]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1687;
      end

       1687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[759] = heapMem[localMem[758]*6 + localMem[757]];
              updateArrayLength(2, 0, 0);
              ip = 1688;
      end

       1688 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[759] != localMem[727] ? 1707 : 1689;
      end

       1689 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[760] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1690;
      end

       1690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[761] = heapMem[localMem[760]*6 + localMem[732]];
              updateArrayLength(2, 0, 0);
              ip = 1691;
      end

       1691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[762] = heapMem[localMem[734]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1692;
      end

       1692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[762]*6 + localMem[757]] = localMem[761];
              updateArrayLength(1, localMem[762], localMem[757]);
              ip = 1693;
      end

       1693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[763] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1694;
      end

       1694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[764] = heapMem[localMem[763]*6 + localMem[732]];
              updateArrayLength(2, 0, 0);
              ip = 1695;
      end

       1695 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[765] = heapMem[localMem[734]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1696;
      end

       1696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[765]*6 + localMem[757]] = localMem[764];
              updateArrayLength(1, localMem[765], localMem[757]);
              ip = 1697;
      end

       1697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[766] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1698;
      end

       1698 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[766]] = localMem[732];
              ip = 1699;
      end

       1699 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[767] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1700;
      end

       1700 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[767]] = localMem[732];
              ip = 1701;
      end

       1701 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[768] = localMem[757] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1702;
      end

       1702 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[734]*6 + 0] = localMem[768];
              updateArrayLength(1, localMem[734], 0);
              ip = 1703;
      end

       1703 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[769] = heapMem[localMem[734]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1704;
      end

       1704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[769]*6 + localMem[768]] = localMem[735];
              updateArrayLength(1, localMem[769], localMem[768]);
              ip = 1705;
      end

       1705 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1845;
      end

       1706 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1729;
      end

       1707 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1708;
      end

       1708 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 1709;
      end

       1709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[770] = heapMem[localMem[734]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1710;
      end

       1710 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[771] = 0; k = arraySizes[localMem[770]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[770] * NArea + i] == localMem[727]) localMem[771] = i + 1;
              end
              ip = 1711;
      end

       1711 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[771] = localMem[771] - 1;
              updateArrayLength(2, 0, 0);
              ip = 1712;
      end

       1712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[772] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1713;
      end

       1713 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[773] = heapMem[localMem[772]*6 + localMem[732]];
              updateArrayLength(2, 0, 0);
              ip = 1714;
      end

       1714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[774] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1715;
      end

       1715 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[775] = heapMem[localMem[774]*6 + localMem[732]];
              updateArrayLength(2, 0, 0);
              ip = 1716;
      end

       1716 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[776] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1717;
      end

       1717 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[776]] = localMem[732];
              ip = 1718;
      end

       1718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[777] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1719;
      end

       1719 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[777]] = localMem[732];
              ip = 1720;
      end

       1720 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[778] = heapMem[localMem[734]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1721;
      end

       1721 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[778] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[771], localMem[778], arraySizes[localMem[778]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[771] && i <= arraySizes[localMem[778]]) begin
                  heapMem[NArea * localMem[778] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[778] + localMem[771]] = localMem[773];                                    // Insert new value
              arraySizes[localMem[778]] = arraySizes[localMem[778]] + 1;                              // Increase array size
              ip = 1722;
      end

       1722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[779] = heapMem[localMem[734]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1723;
      end

       1723 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[779] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[771], localMem[779], arraySizes[localMem[779]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[771] && i <= arraySizes[localMem[779]]) begin
                  heapMem[NArea * localMem[779] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[779] + localMem[771]] = localMem[775];                                    // Insert new value
              arraySizes[localMem[779]] = arraySizes[localMem[779]] + 1;                              // Increase array size
              ip = 1724;
      end

       1724 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[780] = heapMem[localMem[734]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1725;
      end

       1725 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[781] = localMem[771] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1726;
      end

       1726 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[780] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[781], localMem[780], arraySizes[localMem[780]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[781] && i <= arraySizes[localMem[780]]) begin
                  heapMem[NArea * localMem[780] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[780] + localMem[781]] = localMem[735];                                    // Insert new value
              arraySizes[localMem[780]] = arraySizes[localMem[780]] + 1;                              // Increase array size
              ip = 1727;
      end

       1727 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[734]*6 + 0] = heapMem[localMem[734]*6 + 0] + 1;
              updateArrayLength(1, localMem[734], 0);
              ip = 1728;
      end

       1728 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1845;
      end

       1729 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1730;
      end

       1730 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1731;
      end

       1731 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[782] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[782] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[782]] = 0;
              ip = 1732;
      end

       1732 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 0] = localMem[732];
              updateArrayLength(1, localMem[782], 0);
              ip = 1733;
      end

       1733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 2] = 0;
              updateArrayLength(1, localMem[782], 2);
              ip = 1734;
      end

       1734 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[783] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[783] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[783]] = 0;
              ip = 1735;
      end

       1735 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 4] = localMem[783];
              updateArrayLength(1, localMem[782], 4);
              ip = 1736;
      end

       1736 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[784] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[784] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[784]] = 0;
              ip = 1737;
      end

       1737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 5] = localMem[784];
              updateArrayLength(1, localMem[782], 5);
              ip = 1738;
      end

       1738 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 6] = 0;
              updateArrayLength(1, localMem[782], 6);
              ip = 1739;
      end

       1739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 3] = localMem[730];
              updateArrayLength(1, localMem[782], 3);
              ip = 1740;
      end

       1740 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[730]*6 + 1] = heapMem[localMem[730]*6 + 1] + 1;
              updateArrayLength(1, localMem[730], 1);
              ip = 1741;
      end

       1741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 1] = heapMem[localMem[730]*6 + 1];
              updateArrayLength(1, localMem[782], 1);
              ip = 1742;
      end

       1742 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[785] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[785] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[785]] = 0;
              ip = 1743;
      end

       1743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 0] = localMem[732];
              updateArrayLength(1, localMem[785], 0);
              ip = 1744;
      end

       1744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 2] = 0;
              updateArrayLength(1, localMem[785], 2);
              ip = 1745;
      end

       1745 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[786] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[786] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[786]] = 0;
              ip = 1746;
      end

       1746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 4] = localMem[786];
              updateArrayLength(1, localMem[785], 4);
              ip = 1747;
      end

       1747 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[787] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[787] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[787]] = 0;
              ip = 1748;
      end

       1748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 5] = localMem[787];
              updateArrayLength(1, localMem[785], 5);
              ip = 1749;
      end

       1749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 6] = 0;
              updateArrayLength(1, localMem[785], 6);
              ip = 1750;
      end

       1750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 3] = localMem[730];
              updateArrayLength(1, localMem[785], 3);
              ip = 1751;
      end

       1751 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[730]*6 + 1] = heapMem[localMem[730]*6 + 1] + 1;
              updateArrayLength(1, localMem[730], 1);
              ip = 1752;
      end

       1752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 1] = heapMem[localMem[730]*6 + 1];
              updateArrayLength(1, localMem[785], 1);
              ip = 1753;
      end

       1753 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[788] = !heapMem[localMem[727]*6 + 6];
              ip = 1754;
      end

       1754 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[788] != 0 ? 1806 : 1755;
      end

       1755 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[789] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[789] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[789]] = 0;
              ip = 1756;
      end

       1756 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 6] = localMem[789];
              updateArrayLength(1, localMem[782], 6);
              ip = 1757;
      end

       1757 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[790] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[790] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[790]] = 0;
              ip = 1758;
      end

       1758 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 6] = localMem[790];
              updateArrayLength(1, localMem[785], 6);
              ip = 1759;
      end

       1759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[791] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1760;
      end

       1760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[792] = heapMem[localMem[782]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1761;
      end

       1761 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[792] + 0 + i] = heapMem[NArea * localMem[791] + 0 + i];
                  updateArrayLength(1, localMem[792], 0 + i);
                end
              end
              ip = 1762;
      end

       1762 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[793] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1763;
      end

       1763 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[794] = heapMem[localMem[782]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1764;
      end

       1764 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[794] + 0 + i] = heapMem[NArea * localMem[793] + 0 + i];
                  updateArrayLength(1, localMem[794], 0 + i);
                end
              end
              ip = 1765;
      end

       1765 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[795] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1766;
      end

       1766 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[796] = heapMem[localMem[782]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1767;
      end

       1767 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[797] = localMem[732] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1768;
      end

       1768 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[797]) begin
                  heapMem[NArea * localMem[796] + 0 + i] = heapMem[NArea * localMem[795] + 0 + i];
                  updateArrayLength(1, localMem[796], 0 + i);
                end
              end
              ip = 1769;
      end

       1769 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[798] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1770;
      end

       1770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[799] = heapMem[localMem[785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1771;
      end

       1771 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[799] + 0 + i] = heapMem[NArea * localMem[798] + localMem[733] + i];
                  updateArrayLength(1, localMem[799], 0 + i);
                end
              end
              ip = 1772;
      end

       1772 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[800] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1773;
      end

       1773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[801] = heapMem[localMem[785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1774;
      end

       1774 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[801] + 0 + i] = heapMem[NArea * localMem[800] + localMem[733] + i];
                  updateArrayLength(1, localMem[801], 0 + i);
                end
              end
              ip = 1775;
      end

       1775 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[802] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1776;
      end

       1776 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[803] = heapMem[localMem[785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1777;
      end

       1777 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[804] = localMem[732] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1778;
      end

       1778 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[804]) begin
                  heapMem[NArea * localMem[803] + 0 + i] = heapMem[NArea * localMem[802] + localMem[733] + i];
                  updateArrayLength(1, localMem[803], 0 + i);
                end
              end
              ip = 1779;
      end

       1779 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[805] = heapMem[localMem[782]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1780;
      end

       1780 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[806] = localMem[805] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1781;
      end

       1781 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[807] = heapMem[localMem[782]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1782;
      end

       1782 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1783;
      end

       1783 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[808] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1784;
      end

       1784 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1785;
      end

       1785 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[808] >= localMem[806] ? 1791 : 1786;
      end

       1786 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[809] = heapMem[localMem[807]*6 + localMem[808]];
              updateArrayLength(2, 0, 0);
              ip = 1787;
      end

       1787 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[809]*6 + 2] = localMem[782];
              updateArrayLength(1, localMem[809], 2);
              ip = 1788;
      end

       1788 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1789;
      end

       1789 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[808] = localMem[808] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1790;
      end

       1790 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1784;
      end

       1791 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1792;
      end

       1792 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[810] = heapMem[localMem[785]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1793;
      end

       1793 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[811] = localMem[810] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1794;
      end

       1794 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[812] = heapMem[localMem[785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1795;
      end

       1795 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1796;
      end

       1796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[813] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1797;
      end

       1797 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1798;
      end

       1798 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[813] >= localMem[811] ? 1804 : 1799;
      end

       1799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[814] = heapMem[localMem[812]*6 + localMem[813]];
              updateArrayLength(2, 0, 0);
              ip = 1800;
      end

       1800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[814]*6 + 2] = localMem[785];
              updateArrayLength(1, localMem[814], 2);
              ip = 1801;
      end

       1801 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1802;
      end

       1802 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[813] = localMem[813] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1803;
      end

       1803 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1797;
      end

       1804 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1805;
      end

       1805 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1821;
      end

       1806 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1807;
      end

       1807 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[815] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[815] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[815]] = 0;
              ip = 1808;
      end

       1808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[727]*6 + 6] = localMem[815];
              updateArrayLength(1, localMem[727], 6);
              ip = 1809;
      end

       1809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[816] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1810;
      end

       1810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[817] = heapMem[localMem[782]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1811;
      end

       1811 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[817] + 0 + i] = heapMem[NArea * localMem[816] + 0 + i];
                  updateArrayLength(1, localMem[817], 0 + i);
                end
              end
              ip = 1812;
      end

       1812 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[818] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1813;
      end

       1813 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[819] = heapMem[localMem[782]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1814;
      end

       1814 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[819] + 0 + i] = heapMem[NArea * localMem[818] + 0 + i];
                  updateArrayLength(1, localMem[819], 0 + i);
                end
              end
              ip = 1815;
      end

       1815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[820] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1816;
      end

       1816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[821] = heapMem[localMem[785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1817;
      end

       1817 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[821] + 0 + i] = heapMem[NArea * localMem[820] + localMem[733] + i];
                  updateArrayLength(1, localMem[821], 0 + i);
                end
              end
              ip = 1818;
      end

       1818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[822] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1819;
      end

       1819 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[823] = heapMem[localMem[785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1820;
      end

       1820 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[732]) begin
                  heapMem[NArea * localMem[823] + 0 + i] = heapMem[NArea * localMem[822] + localMem[733] + i];
                  updateArrayLength(1, localMem[823], 0 + i);
                end
              end
              ip = 1821;
      end

       1821 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1822;
      end

       1822 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[782]*6 + 2] = localMem[727];
              updateArrayLength(1, localMem[782], 2);
              ip = 1823;
      end

       1823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[785]*6 + 2] = localMem[727];
              updateArrayLength(1, localMem[785], 2);
              ip = 1824;
      end

       1824 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[824] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1825;
      end

       1825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[825] = heapMem[localMem[824]*6 + localMem[732]];
              updateArrayLength(2, 0, 0);
              ip = 1826;
      end

       1826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[826] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1827;
      end

       1827 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[827] = heapMem[localMem[826]*6 + localMem[732]];
              updateArrayLength(2, 0, 0);
              ip = 1828;
      end

       1828 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[828] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1829;
      end

       1829 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[828]*6 + 0] = localMem[825];
              updateArrayLength(1, localMem[828], 0);
              ip = 1830;
      end

       1830 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[829] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1831;
      end

       1831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[829]*6 + 0] = localMem[827];
              updateArrayLength(1, localMem[829], 0);
              ip = 1832;
      end

       1832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[830] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1833;
      end

       1833 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[830]*6 + 0] = localMem[782];
              updateArrayLength(1, localMem[830], 0);
              ip = 1834;
      end

       1834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[831] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1835;
      end

       1835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[831]*6 + 1] = localMem[785];
              updateArrayLength(1, localMem[831], 1);
              ip = 1836;
      end

       1836 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[727]*6 + 0] = 1;
              updateArrayLength(1, localMem[727], 0);
              ip = 1837;
      end

       1837 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[832] = heapMem[localMem[727]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1838;
      end

       1838 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[832]] = 1;
              ip = 1839;
      end

       1839 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[833] = heapMem[localMem[727]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1840;
      end

       1840 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[833]] = 1;
              ip = 1841;
      end

       1841 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[834] = heapMem[localMem[727]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1842;
      end

       1842 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[834]] = 2;
              ip = 1843;
      end

       1843 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1845;
      end

       1844 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1850;
      end

       1845 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1846;
      end

       1846 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[728] = 1;
              updateArrayLength(2, 0, 0);
              ip = 1847;
      end

       1847 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1850;
      end

       1848 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1849;
      end

       1849 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[728] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1850;
      end

       1850 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1851;
      end

       1851 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[728] != 0 ? 1853 : 1852;
      end

       1852 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[499] = localMem[727];
              updateArrayLength(2, 0, 0);
              ip = 1853;
      end

       1853 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1854;
      end

       1854 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1855;
      end

       1855 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[607] = localMem[607] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1856;
      end

       1856 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1358;
      end

       1857 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1858;
      end

       1858 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
            ip = 1859;
      end

       1859 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1860;
      end

       1860 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1861;
      end

       1861 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1862;
      end

       1862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[835] = heapMem[localMem[476]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1863;
      end

       1863 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[836] = heapMem[localMem[476]*6 + 1];
              updateArrayLength(2, 0, 0);
              ip = 1864;
      end

       1864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[837] = heapMem[localMem[476]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1865;
      end

       1865 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[836] != 1 ? 1869 : 1866;
      end

       1866 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[838] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1867;
      end

       1867 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[838]*6 + localMem[837]] = 22;
              updateArrayLength(1, localMem[838], localMem[837]);
              ip = 1868;
      end

       1868 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2115;
      end

       1869 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1870;
      end

       1870 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[836] != 2 ? 1878 : 1871;
      end

       1871 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[839] = localMem[837] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1872;
      end

       1872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[840] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1873;
      end

       1873 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[840] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[839], localMem[840], arraySizes[localMem[840]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[839] && i <= arraySizes[localMem[840]]) begin
                  heapMem[NArea * localMem[840] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[840] + localMem[839]] = 2;                                    // Insert new value
              arraySizes[localMem[840]] = arraySizes[localMem[840]] + 1;                              // Increase array size
              ip = 1874;
      end

       1874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[841] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1875;
      end

       1875 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[841] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[839], localMem[841], arraySizes[localMem[841]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[839] && i <= arraySizes[localMem[841]]) begin
                  heapMem[NArea * localMem[841] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[841] + localMem[839]] = 22;                                    // Insert new value
              arraySizes[localMem[841]] = arraySizes[localMem[841]] + 1;                              // Increase array size
              ip = 1876;
      end

       1876 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[835]*6 + 0] = heapMem[localMem[835]*6 + 0] + 1;
              updateArrayLength(1, localMem[835], 0);
              ip = 1877;
      end

       1877 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1884;
      end

       1878 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1879;
      end

       1879 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[842] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1880;
      end

       1880 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[842] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[837], localMem[842], arraySizes[localMem[842]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[837] && i <= arraySizes[localMem[842]]) begin
                  heapMem[NArea * localMem[842] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[842] + localMem[837]] = 2;                                    // Insert new value
              arraySizes[localMem[842]] = arraySizes[localMem[842]] + 1;                              // Increase array size
              ip = 1881;
      end

       1881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[843] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1882;
      end

       1882 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[843] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[837], localMem[843], arraySizes[localMem[843]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[837] && i <= arraySizes[localMem[843]]) begin
                  heapMem[NArea * localMem[843] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[843] + localMem[837]] = 22;                                    // Insert new value
              arraySizes[localMem[843]] = arraySizes[localMem[843]] + 1;                              // Increase array size
              ip = 1883;
      end

       1883 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[835]*6 + 0] = heapMem[localMem[835]*6 + 0] + 1;
              updateArrayLength(1, localMem[835], 0);
              ip = 1884;
      end

       1884 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1885;
      end

       1885 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 1886;
      end

       1886 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1887;
      end

       1887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[845] = heapMem[localMem[835]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1888;
      end

       1888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[846] = heapMem[localMem[835]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1889;
      end

       1889 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[847] = heapMem[localMem[846]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1890;
      end

       1890 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[845] <  localMem[847] ? 2110 : 1891;
      end

       1891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[848] = localMem[847];
              updateArrayLength(2, 0, 0);
              ip = 1892;
      end

       1892 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[848] = localMem[848] >> 1;
              ip = 1893;
      end

       1893 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[849] = localMem[848] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1894;
      end

       1894 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[850] = heapMem[localMem[835]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1895;
      end

       1895 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[850] == 0 ? 1992 : 1896;
      end

       1896 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[851] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[851] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[851]] = 0;
              ip = 1897;
      end

       1897 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 0] = localMem[848];
              updateArrayLength(1, localMem[851], 0);
              ip = 1898;
      end

       1898 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 2] = 0;
              updateArrayLength(1, localMem[851], 2);
              ip = 1899;
      end

       1899 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[852] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[852] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[852]] = 0;
              ip = 1900;
      end

       1900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 4] = localMem[852];
              updateArrayLength(1, localMem[851], 4);
              ip = 1901;
      end

       1901 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[853] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[853] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[853]] = 0;
              ip = 1902;
      end

       1902 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 5] = localMem[853];
              updateArrayLength(1, localMem[851], 5);
              ip = 1903;
      end

       1903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 6] = 0;
              updateArrayLength(1, localMem[851], 6);
              ip = 1904;
      end

       1904 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 3] = localMem[846];
              updateArrayLength(1, localMem[851], 3);
              ip = 1905;
      end

       1905 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[846]*6 + 1] = heapMem[localMem[846]*6 + 1] + 1;
              updateArrayLength(1, localMem[846], 1);
              ip = 1906;
      end

       1906 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 1] = heapMem[localMem[846]*6 + 1];
              updateArrayLength(1, localMem[851], 1);
              ip = 1907;
      end

       1907 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[854] = !heapMem[localMem[835]*6 + 6];
              ip = 1908;
      end

       1908 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[854] != 0 ? 1937 : 1909;
      end

       1909 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[855] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[855] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[855]] = 0;
              ip = 1910;
      end

       1910 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 6] = localMem[855];
              updateArrayLength(1, localMem[851], 6);
              ip = 1911;
      end

       1911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[856] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1912;
      end

       1912 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[857] = heapMem[localMem[851]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1913;
      end

       1913 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[857] + 0 + i] = heapMem[NArea * localMem[856] + localMem[849] + i];
                  updateArrayLength(1, localMem[857], 0 + i);
                end
              end
              ip = 1914;
      end

       1914 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[858] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1915;
      end

       1915 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[859] = heapMem[localMem[851]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1916;
      end

       1916 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[859] + 0 + i] = heapMem[NArea * localMem[858] + localMem[849] + i];
                  updateArrayLength(1, localMem[859], 0 + i);
                end
              end
              ip = 1917;
      end

       1917 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[860] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1918;
      end

       1918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[861] = heapMem[localMem[851]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1919;
      end

       1919 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[862] = localMem[848] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1920;
      end

       1920 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[862]) begin
                  heapMem[NArea * localMem[861] + 0 + i] = heapMem[NArea * localMem[860] + localMem[849] + i];
                  updateArrayLength(1, localMem[861], 0 + i);
                end
              end
              ip = 1921;
      end

       1921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[863] = heapMem[localMem[851]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1922;
      end

       1922 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[864] = localMem[863] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1923;
      end

       1923 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[865] = heapMem[localMem[851]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1924;
      end

       1924 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1925;
      end

       1925 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[866] = 0;
              updateArrayLength(2, 0, 0);
              ip = 1926;
      end

       1926 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1927;
      end

       1927 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[866] >= localMem[864] ? 1933 : 1928;
      end

       1928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[867] = heapMem[localMem[865]*6 + localMem[866]];
              updateArrayLength(2, 0, 0);
              ip = 1929;
      end

       1929 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[867]*6 + 2] = localMem[851];
              updateArrayLength(1, localMem[867], 2);
              ip = 1930;
      end

       1930 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1931;
      end

       1931 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[866] = localMem[866] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1932;
      end

       1932 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1926;
      end

       1933 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1934;
      end

       1934 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[868] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1935;
      end

       1935 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[868]] = localMem[849];
              ip = 1936;
      end

       1936 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1944;
      end

       1937 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1938;
      end

       1938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[869] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1939;
      end

       1939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[870] = heapMem[localMem[851]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1940;
      end

       1940 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[870] + 0 + i] = heapMem[NArea * localMem[869] + localMem[849] + i];
                  updateArrayLength(1, localMem[870], 0 + i);
                end
              end
              ip = 1941;
      end

       1941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[871] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1942;
      end

       1942 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[872] = heapMem[localMem[851]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1943;
      end

       1943 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[872] + 0 + i] = heapMem[NArea * localMem[871] + localMem[849] + i];
                  updateArrayLength(1, localMem[872], 0 + i);
                end
              end
              ip = 1944;
      end

       1944 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1945;
      end

       1945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[835]*6 + 0] = localMem[848];
              updateArrayLength(1, localMem[835], 0);
              ip = 1946;
      end

       1946 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[851]*6 + 2] = localMem[850];
              updateArrayLength(1, localMem[851], 2);
              ip = 1947;
      end

       1947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[873] = heapMem[localMem[850]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1948;
      end

       1948 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[874] = heapMem[localMem[850]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1949;
      end

       1949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[875] = heapMem[localMem[874]*6 + localMem[873]];
              updateArrayLength(2, 0, 0);
              ip = 1950;
      end

       1950 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[875] != localMem[835] ? 1969 : 1951;
      end

       1951 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[876] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1952;
      end

       1952 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[877] = heapMem[localMem[876]*6 + localMem[848]];
              updateArrayLength(2, 0, 0);
              ip = 1953;
      end

       1953 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[878] = heapMem[localMem[850]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1954;
      end

       1954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[878]*6 + localMem[873]] = localMem[877];
              updateArrayLength(1, localMem[878], localMem[873]);
              ip = 1955;
      end

       1955 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[879] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1956;
      end

       1956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[880] = heapMem[localMem[879]*6 + localMem[848]];
              updateArrayLength(2, 0, 0);
              ip = 1957;
      end

       1957 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[881] = heapMem[localMem[850]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1958;
      end

       1958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[881]*6 + localMem[873]] = localMem[880];
              updateArrayLength(1, localMem[881], localMem[873]);
              ip = 1959;
      end

       1959 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[882] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1960;
      end

       1960 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[882]] = localMem[848];
              ip = 1961;
      end

       1961 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[883] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1962;
      end

       1962 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[883]] = localMem[848];
              ip = 1963;
      end

       1963 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[884] = localMem[873] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1964;
      end

       1964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[850]*6 + 0] = localMem[884];
              updateArrayLength(1, localMem[850], 0);
              ip = 1965;
      end

       1965 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[885] = heapMem[localMem[850]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1966;
      end

       1966 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[885]*6 + localMem[884]] = localMem[851];
              updateArrayLength(1, localMem[885], localMem[884]);
              ip = 1967;
      end

       1967 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2107;
      end

       1968 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1991;
      end

       1969 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1970;
      end

       1970 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 1971;
      end

       1971 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[886] = heapMem[localMem[850]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1972;
      end

       1972 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[887] = 0; k = arraySizes[localMem[886]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[886] * NArea + i] == localMem[835]) localMem[887] = i + 1;
              end
              ip = 1973;
      end

       1973 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[887] = localMem[887] - 1;
              updateArrayLength(2, 0, 0);
              ip = 1974;
      end

       1974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[888] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1975;
      end

       1975 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[889] = heapMem[localMem[888]*6 + localMem[848]];
              updateArrayLength(2, 0, 0);
              ip = 1976;
      end

       1976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[890] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1977;
      end

       1977 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[891] = heapMem[localMem[890]*6 + localMem[848]];
              updateArrayLength(2, 0, 0);
              ip = 1978;
      end

       1978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[892] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1979;
      end

       1979 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[892]] = localMem[848];
              ip = 1980;
      end

       1980 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[893] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1981;
      end

       1981 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[893]] = localMem[848];
              ip = 1982;
      end

       1982 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[894] = heapMem[localMem[850]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1983;
      end

       1983 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[894] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[887], localMem[894], arraySizes[localMem[894]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[887] && i <= arraySizes[localMem[894]]) begin
                  heapMem[NArea * localMem[894] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[894] + localMem[887]] = localMem[889];                                    // Insert new value
              arraySizes[localMem[894]] = arraySizes[localMem[894]] + 1;                              // Increase array size
              ip = 1984;
      end

       1984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[895] = heapMem[localMem[850]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1985;
      end

       1985 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[895] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[887], localMem[895], arraySizes[localMem[895]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[887] && i <= arraySizes[localMem[895]]) begin
                  heapMem[NArea * localMem[895] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[895] + localMem[887]] = localMem[891];                                    // Insert new value
              arraySizes[localMem[895]] = arraySizes[localMem[895]] + 1;                              // Increase array size
              ip = 1986;
      end

       1986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[896] = heapMem[localMem[850]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 1987;
      end

       1987 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[897] = localMem[887] + 1;
              updateArrayLength(2, 0, 0);
              ip = 1988;
      end

       1988 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[896] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[897], localMem[896], arraySizes[localMem[896]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[897] && i <= arraySizes[localMem[896]]) begin
                  heapMem[NArea * localMem[896] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[896] + localMem[897]] = localMem[851];                                    // Insert new value
              arraySizes[localMem[896]] = arraySizes[localMem[896]] + 1;                              // Increase array size
              ip = 1989;
      end

       1989 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[850]*6 + 0] = heapMem[localMem[850]*6 + 0] + 1;
              updateArrayLength(1, localMem[850], 0);
              ip = 1990;
      end

       1990 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2107;
      end

       1991 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1992;
      end

       1992 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1993;
      end

       1993 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[898] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[898] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[898]] = 0;
              ip = 1994;
      end

       1994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 0] = localMem[848];
              updateArrayLength(1, localMem[898], 0);
              ip = 1995;
      end

       1995 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 2] = 0;
              updateArrayLength(1, localMem[898], 2);
              ip = 1996;
      end

       1996 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[899] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[899] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[899]] = 0;
              ip = 1997;
      end

       1997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 4] = localMem[899];
              updateArrayLength(1, localMem[898], 4);
              ip = 1998;
      end

       1998 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[900] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[900] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[900]] = 0;
              ip = 1999;
      end

       1999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 5] = localMem[900];
              updateArrayLength(1, localMem[898], 5);
              ip = 2000;
      end

       2000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 6] = 0;
              updateArrayLength(1, localMem[898], 6);
              ip = 2001;
      end

       2001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 3] = localMem[846];
              updateArrayLength(1, localMem[898], 3);
              ip = 2002;
      end

       2002 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[846]*6 + 1] = heapMem[localMem[846]*6 + 1] + 1;
              updateArrayLength(1, localMem[846], 1);
              ip = 2003;
      end

       2003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 1] = heapMem[localMem[846]*6 + 1];
              updateArrayLength(1, localMem[898], 1);
              ip = 2004;
      end

       2004 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[901] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[901] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[901]] = 0;
              ip = 2005;
      end

       2005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 0] = localMem[848];
              updateArrayLength(1, localMem[901], 0);
              ip = 2006;
      end

       2006 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 2] = 0;
              updateArrayLength(1, localMem[901], 2);
              ip = 2007;
      end

       2007 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[902] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[902] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[902]] = 0;
              ip = 2008;
      end

       2008 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 4] = localMem[902];
              updateArrayLength(1, localMem[901], 4);
              ip = 2009;
      end

       2009 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[903] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[903] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[903]] = 0;
              ip = 2010;
      end

       2010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 5] = localMem[903];
              updateArrayLength(1, localMem[901], 5);
              ip = 2011;
      end

       2011 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 6] = 0;
              updateArrayLength(1, localMem[901], 6);
              ip = 2012;
      end

       2012 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 3] = localMem[846];
              updateArrayLength(1, localMem[901], 3);
              ip = 2013;
      end

       2013 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[846]*6 + 1] = heapMem[localMem[846]*6 + 1] + 1;
              updateArrayLength(1, localMem[846], 1);
              ip = 2014;
      end

       2014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 1] = heapMem[localMem[846]*6 + 1];
              updateArrayLength(1, localMem[901], 1);
              ip = 2015;
      end

       2015 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[904] = !heapMem[localMem[835]*6 + 6];
              ip = 2016;
      end

       2016 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[904] != 0 ? 2068 : 2017;
      end

       2017 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[905] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[905] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[905]] = 0;
              ip = 2018;
      end

       2018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 6] = localMem[905];
              updateArrayLength(1, localMem[898], 6);
              ip = 2019;
      end

       2019 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[906] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[906] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[906]] = 0;
              ip = 2020;
      end

       2020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 6] = localMem[906];
              updateArrayLength(1, localMem[901], 6);
              ip = 2021;
      end

       2021 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[907] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2022;
      end

       2022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[908] = heapMem[localMem[898]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2023;
      end

       2023 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[908] + 0 + i] = heapMem[NArea * localMem[907] + 0 + i];
                  updateArrayLength(1, localMem[908], 0 + i);
                end
              end
              ip = 2024;
      end

       2024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[909] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2025;
      end

       2025 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[910] = heapMem[localMem[898]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2026;
      end

       2026 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[910] + 0 + i] = heapMem[NArea * localMem[909] + 0 + i];
                  updateArrayLength(1, localMem[910], 0 + i);
                end
              end
              ip = 2027;
      end

       2027 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[911] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2028;
      end

       2028 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[912] = heapMem[localMem[898]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2029;
      end

       2029 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[913] = localMem[848] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2030;
      end

       2030 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[913]) begin
                  heapMem[NArea * localMem[912] + 0 + i] = heapMem[NArea * localMem[911] + 0 + i];
                  updateArrayLength(1, localMem[912], 0 + i);
                end
              end
              ip = 2031;
      end

       2031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[914] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2032;
      end

       2032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[915] = heapMem[localMem[901]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2033;
      end

       2033 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[915] + 0 + i] = heapMem[NArea * localMem[914] + localMem[849] + i];
                  updateArrayLength(1, localMem[915], 0 + i);
                end
              end
              ip = 2034;
      end

       2034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[916] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2035;
      end

       2035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[917] = heapMem[localMem[901]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2036;
      end

       2036 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[917] + 0 + i] = heapMem[NArea * localMem[916] + localMem[849] + i];
                  updateArrayLength(1, localMem[917], 0 + i);
                end
              end
              ip = 2037;
      end

       2037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[918] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2038;
      end

       2038 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[919] = heapMem[localMem[901]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2039;
      end

       2039 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[920] = localMem[848] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2040;
      end

       2040 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[920]) begin
                  heapMem[NArea * localMem[919] + 0 + i] = heapMem[NArea * localMem[918] + localMem[849] + i];
                  updateArrayLength(1, localMem[919], 0 + i);
                end
              end
              ip = 2041;
      end

       2041 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[921] = heapMem[localMem[898]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2042;
      end

       2042 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[922] = localMem[921] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2043;
      end

       2043 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[923] = heapMem[localMem[898]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2044;
      end

       2044 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2045;
      end

       2045 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[924] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2046;
      end

       2046 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2047;
      end

       2047 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[924] >= localMem[922] ? 2053 : 2048;
      end

       2048 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[925] = heapMem[localMem[923]*6 + localMem[924]];
              updateArrayLength(2, 0, 0);
              ip = 2049;
      end

       2049 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[925]*6 + 2] = localMem[898];
              updateArrayLength(1, localMem[925], 2);
              ip = 2050;
      end

       2050 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2051;
      end

       2051 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[924] = localMem[924] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2052;
      end

       2052 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2046;
      end

       2053 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2054;
      end

       2054 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[926] = heapMem[localMem[901]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2055;
      end

       2055 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[927] = localMem[926] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2056;
      end

       2056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[928] = heapMem[localMem[901]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2057;
      end

       2057 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2058;
      end

       2058 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[929] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2059;
      end

       2059 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2060;
      end

       2060 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[929] >= localMem[927] ? 2066 : 2061;
      end

       2061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[930] = heapMem[localMem[928]*6 + localMem[929]];
              updateArrayLength(2, 0, 0);
              ip = 2062;
      end

       2062 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[930]*6 + 2] = localMem[901];
              updateArrayLength(1, localMem[930], 2);
              ip = 2063;
      end

       2063 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2064;
      end

       2064 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[929] = localMem[929] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2065;
      end

       2065 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2059;
      end

       2066 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2067;
      end

       2067 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2083;
      end

       2068 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2069;
      end

       2069 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[931] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[931] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[931]] = 0;
              ip = 2070;
      end

       2070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[835]*6 + 6] = localMem[931];
              updateArrayLength(1, localMem[835], 6);
              ip = 2071;
      end

       2071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[932] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2072;
      end

       2072 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[933] = heapMem[localMem[898]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2073;
      end

       2073 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[933] + 0 + i] = heapMem[NArea * localMem[932] + 0 + i];
                  updateArrayLength(1, localMem[933], 0 + i);
                end
              end
              ip = 2074;
      end

       2074 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[934] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2075;
      end

       2075 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[935] = heapMem[localMem[898]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2076;
      end

       2076 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[935] + 0 + i] = heapMem[NArea * localMem[934] + 0 + i];
                  updateArrayLength(1, localMem[935], 0 + i);
                end
              end
              ip = 2077;
      end

       2077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[936] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2078;
      end

       2078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[937] = heapMem[localMem[901]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2079;
      end

       2079 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[937] + 0 + i] = heapMem[NArea * localMem[936] + localMem[849] + i];
                  updateArrayLength(1, localMem[937], 0 + i);
                end
              end
              ip = 2080;
      end

       2080 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[938] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2081;
      end

       2081 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[939] = heapMem[localMem[901]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2082;
      end

       2082 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[848]) begin
                  heapMem[NArea * localMem[939] + 0 + i] = heapMem[NArea * localMem[938] + localMem[849] + i];
                  updateArrayLength(1, localMem[939], 0 + i);
                end
              end
              ip = 2083;
      end

       2083 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2084;
      end

       2084 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[898]*6 + 2] = localMem[835];
              updateArrayLength(1, localMem[898], 2);
              ip = 2085;
      end

       2085 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[901]*6 + 2] = localMem[835];
              updateArrayLength(1, localMem[901], 2);
              ip = 2086;
      end

       2086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[940] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2087;
      end

       2087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[941] = heapMem[localMem[940]*6 + localMem[848]];
              updateArrayLength(2, 0, 0);
              ip = 2088;
      end

       2088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[942] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2089;
      end

       2089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[943] = heapMem[localMem[942]*6 + localMem[848]];
              updateArrayLength(2, 0, 0);
              ip = 2090;
      end

       2090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[944] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2091;
      end

       2091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[944]*6 + 0] = localMem[941];
              updateArrayLength(1, localMem[944], 0);
              ip = 2092;
      end

       2092 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[945] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2093;
      end

       2093 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[945]*6 + 0] = localMem[943];
              updateArrayLength(1, localMem[945], 0);
              ip = 2094;
      end

       2094 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[946] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2095;
      end

       2095 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[946]*6 + 0] = localMem[898];
              updateArrayLength(1, localMem[946], 0);
              ip = 2096;
      end

       2096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[947] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2097;
      end

       2097 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[947]*6 + 1] = localMem[901];
              updateArrayLength(1, localMem[947], 1);
              ip = 2098;
      end

       2098 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[835]*6 + 0] = 1;
              updateArrayLength(1, localMem[835], 0);
              ip = 2099;
      end

       2099 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[948] = heapMem[localMem[835]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2100;
      end

       2100 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[948]] = 1;
              ip = 2101;
      end

       2101 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[949] = heapMem[localMem[835]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2102;
      end

       2102 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[949]] = 1;
              ip = 2103;
      end

       2103 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[950] = heapMem[localMem[835]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2104;
      end

       2104 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[950]] = 2;
              ip = 2105;
      end

       2105 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2107;
      end

       2106 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2112;
      end

       2107 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2108;
      end

       2108 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[844] = 1;
              updateArrayLength(2, 0, 0);
              ip = 2109;
      end

       2109 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2112;
      end

       2110 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2111;
      end

       2111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[844] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2112;
      end

       2112 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2113;
      end

       2113 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2114;
      end

       2114 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2115;
      end

       2115 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2116;
      end

       2116 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[476]] = 0;
              freedArrays[freedArraysTop] = localMem[476];
              freedArraysTop = freedArraysTop + 1;
              ip = 2117;
      end

       2117 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[951] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[951] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[951]] = 0;
              ip = 2118;
      end

       2118 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2119;
      end

       2119 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[952] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2120;
      end

       2120 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[952] != 0 ? 2143 : 2121;
      end

       2121 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[953] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[953] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[953]] = 0;
              ip = 2122;
      end

       2122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 0] = 1;
              updateArrayLength(1, localMem[953], 0);
              ip = 2123;
      end

       2123 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 2] = 0;
              updateArrayLength(1, localMem[953], 2);
              ip = 2124;
      end

       2124 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[954] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[954] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[954]] = 0;
              ip = 2125;
      end

       2125 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 4] = localMem[954];
              updateArrayLength(1, localMem[953], 4);
              ip = 2126;
      end

       2126 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[955] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[955] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[955]] = 0;
              ip = 2127;
      end

       2127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 5] = localMem[955];
              updateArrayLength(1, localMem[953], 5);
              ip = 2128;
      end

       2128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 6] = 0;
              updateArrayLength(1, localMem[953], 6);
              ip = 2129;
      end

       2129 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 3] = localMem[0];
              updateArrayLength(1, localMem[953], 3);
              ip = 2130;
      end

       2130 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = heapMem[localMem[0]*6 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 2131;
      end

       2131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[953]*6 + 1] = heapMem[localMem[0]*6 + 1];
              updateArrayLength(1, localMem[953], 1);
              ip = 2132;
      end

       2132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[956] = heapMem[localMem[953]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2133;
      end

       2133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[956]*6 + 0] = 3;
              updateArrayLength(1, localMem[956], 0);
              ip = 2134;
      end

       2134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[957] = heapMem[localMem[953]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2135;
      end

       2135 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[957]*6 + 0] = 33;
              updateArrayLength(1, localMem[957], 0);
              ip = 2136;
      end

       2136 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 2137;
      end

       2137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = localMem[953];
              updateArrayLength(1, localMem[0], 3);
              ip = 2138;
      end

       2138 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[958] = heapMem[localMem[953]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2139;
      end

       2139 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[958]] = 1;
              ip = 2140;
      end

       2140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[959] = heapMem[localMem[953]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2141;
      end

       2141 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[959]] = 1;
              ip = 2142;
      end

       2142 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3171;
      end

       2143 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2144;
      end

       2144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[960] = heapMem[localMem[952]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2145;
      end

       2145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[961] = heapMem[localMem[0]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2146;
      end

       2146 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[960] >= localMem[961] ? 2182 : 2147;
      end

       2147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[962] = heapMem[localMem[952]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2148;
      end

       2148 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[962] != 0 ? 2181 : 2149;
      end

       2149 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[963] = !heapMem[localMem[952]*6 + 6];
              ip = 2150;
      end

       2150 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[963] == 0 ? 2180 : 2151;
      end

       2151 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[964] = heapMem[localMem[952]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2152;
      end

       2152 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[965] = 0; k = arraySizes[localMem[964]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[964] * NArea + i] == 3) localMem[965] = i + 1;
              end
              ip = 2153;
      end

       2153 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[965] == 0 ? 2158 : 2154;
      end

       2154 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[965] = localMem[965] - 1;
              updateArrayLength(2, 0, 0);
              ip = 2155;
      end

       2155 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[966] = heapMem[localMem[952]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2156;
      end

       2156 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[966]*6 + localMem[965]] = 33;
              updateArrayLength(1, localMem[966], localMem[965]);
              ip = 2157;
      end

       2157 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3171;
      end

       2158 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2159;
      end

       2159 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[964]] = localMem[960];
              ip = 2160;
      end

       2160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[967] = heapMem[localMem[952]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2161;
      end

       2161 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[967]] = localMem[960];
              ip = 2162;
      end

       2162 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[964]];
//$display("AAAAA k=%d  source2=%d", k, 3);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[964] * NArea + i]);
                if (i < k && heapMem[localMem[964] * NArea + i] > 3) j = j + 1;
              end
              localMem[968] = j;
              ip = 2163;
      end

       2163 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[968] != 0 ? 2171 : 2164;
      end

       2164 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[969] = heapMem[localMem[952]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2165;
      end

       2165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[969]*6 + localMem[960]] = 3;
              updateArrayLength(1, localMem[969], localMem[960]);
              ip = 2166;
      end

       2166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[970] = heapMem[localMem[952]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2167;
      end

       2167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[970]*6 + localMem[960]] = 33;
              updateArrayLength(1, localMem[970], localMem[960]);
              ip = 2168;
      end

       2168 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[952]*6 + 0] = localMem[960] + 1;
              updateArrayLength(1, localMem[952], 0);
              ip = 2169;
      end

       2169 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 2170;
      end

       2170 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3171;
      end

       2171 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2172;
      end

       2172 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[964]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[964] * NArea + i] < 3) j = j + 1;
              end
              localMem[971] = j;
              ip = 2173;
      end

       2173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[972] = heapMem[localMem[952]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2174;
      end

       2174 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[972] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[971], localMem[972], arraySizes[localMem[972]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[971] && i <= arraySizes[localMem[972]]) begin
                  heapMem[NArea * localMem[972] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[972] + localMem[971]] = 3;                                    // Insert new value
              arraySizes[localMem[972]] = arraySizes[localMem[972]] + 1;                              // Increase array size
              ip = 2175;
      end

       2175 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[973] = heapMem[localMem[952]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2176;
      end

       2176 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[973] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[971], localMem[973], arraySizes[localMem[973]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[971] && i <= arraySizes[localMem[973]]) begin
                  heapMem[NArea * localMem[973] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[973] + localMem[971]] = 33;                                    // Insert new value
              arraySizes[localMem[973]] = arraySizes[localMem[973]] + 1;                              // Increase array size
              ip = 2177;
      end

       2177 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[952]*6 + 0] = heapMem[localMem[952]*6 + 0] + 1;
              updateArrayLength(1, localMem[952], 0);
              ip = 2178;
      end

       2178 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 2179;
      end

       2179 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3171;
      end

       2180 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2181;
      end

       2181 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2182;
      end

       2182 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2183;
      end

       2183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[974] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2184;
      end

       2184 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2185;
      end

       2185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[976] = heapMem[localMem[974]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2186;
      end

       2186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[977] = heapMem[localMem[974]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2187;
      end

       2187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[978] = heapMem[localMem[977]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2188;
      end

       2188 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[976] <  localMem[978] ? 2408 : 2189;
      end

       2189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[979] = localMem[978];
              updateArrayLength(2, 0, 0);
              ip = 2190;
      end

       2190 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[979] = localMem[979] >> 1;
              ip = 2191;
      end

       2191 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[980] = localMem[979] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2192;
      end

       2192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[981] = heapMem[localMem[974]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2193;
      end

       2193 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[981] == 0 ? 2290 : 2194;
      end

       2194 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[982] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[982] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[982]] = 0;
              ip = 2195;
      end

       2195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 0] = localMem[979];
              updateArrayLength(1, localMem[982], 0);
              ip = 2196;
      end

       2196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 2] = 0;
              updateArrayLength(1, localMem[982], 2);
              ip = 2197;
      end

       2197 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[983] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[983] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[983]] = 0;
              ip = 2198;
      end

       2198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 4] = localMem[983];
              updateArrayLength(1, localMem[982], 4);
              ip = 2199;
      end

       2199 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[984] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[984] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[984]] = 0;
              ip = 2200;
      end

       2200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 5] = localMem[984];
              updateArrayLength(1, localMem[982], 5);
              ip = 2201;
      end

       2201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 6] = 0;
              updateArrayLength(1, localMem[982], 6);
              ip = 2202;
      end

       2202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 3] = localMem[977];
              updateArrayLength(1, localMem[982], 3);
              ip = 2203;
      end

       2203 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[977]*6 + 1] = heapMem[localMem[977]*6 + 1] + 1;
              updateArrayLength(1, localMem[977], 1);
              ip = 2204;
      end

       2204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 1] = heapMem[localMem[977]*6 + 1];
              updateArrayLength(1, localMem[982], 1);
              ip = 2205;
      end

       2205 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[985] = !heapMem[localMem[974]*6 + 6];
              ip = 2206;
      end

       2206 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[985] != 0 ? 2235 : 2207;
      end

       2207 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[986] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[986] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[986]] = 0;
              ip = 2208;
      end

       2208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 6] = localMem[986];
              updateArrayLength(1, localMem[982], 6);
              ip = 2209;
      end

       2209 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[987] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2210;
      end

       2210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[988] = heapMem[localMem[982]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2211;
      end

       2211 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[988] + 0 + i] = heapMem[NArea * localMem[987] + localMem[980] + i];
                  updateArrayLength(1, localMem[988], 0 + i);
                end
              end
              ip = 2212;
      end

       2212 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[989] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2213;
      end

       2213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[990] = heapMem[localMem[982]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2214;
      end

       2214 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[990] + 0 + i] = heapMem[NArea * localMem[989] + localMem[980] + i];
                  updateArrayLength(1, localMem[990], 0 + i);
                end
              end
              ip = 2215;
      end

       2215 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[991] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2216;
      end

       2216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[992] = heapMem[localMem[982]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2217;
      end

       2217 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[993] = localMem[979] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2218;
      end

       2218 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[993]) begin
                  heapMem[NArea * localMem[992] + 0 + i] = heapMem[NArea * localMem[991] + localMem[980] + i];
                  updateArrayLength(1, localMem[992], 0 + i);
                end
              end
              ip = 2219;
      end

       2219 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[994] = heapMem[localMem[982]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2220;
      end

       2220 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[995] = localMem[994] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2221;
      end

       2221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[996] = heapMem[localMem[982]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2222;
      end

       2222 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2223;
      end

       2223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[997] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2224;
      end

       2224 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2225;
      end

       2225 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[997] >= localMem[995] ? 2231 : 2226;
      end

       2226 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[998] = heapMem[localMem[996]*6 + localMem[997]];
              updateArrayLength(2, 0, 0);
              ip = 2227;
      end

       2227 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[998]*6 + 2] = localMem[982];
              updateArrayLength(1, localMem[998], 2);
              ip = 2228;
      end

       2228 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2229;
      end

       2229 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[997] = localMem[997] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2230;
      end

       2230 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2224;
      end

       2231 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2232;
      end

       2232 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[999] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2233;
      end

       2233 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[999]] = localMem[980];
              ip = 2234;
      end

       2234 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2242;
      end

       2235 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2236;
      end

       2236 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1000] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2237;
      end

       2237 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1001] = heapMem[localMem[982]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2238;
      end

       2238 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1001] + 0 + i] = heapMem[NArea * localMem[1000] + localMem[980] + i];
                  updateArrayLength(1, localMem[1001], 0 + i);
                end
              end
              ip = 2239;
      end

       2239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1002] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2240;
      end

       2240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1003] = heapMem[localMem[982]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2241;
      end

       2241 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1003] + 0 + i] = heapMem[NArea * localMem[1002] + localMem[980] + i];
                  updateArrayLength(1, localMem[1003], 0 + i);
                end
              end
              ip = 2242;
      end

       2242 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2243;
      end

       2243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[974]*6 + 0] = localMem[979];
              updateArrayLength(1, localMem[974], 0);
              ip = 2244;
      end

       2244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[982]*6 + 2] = localMem[981];
              updateArrayLength(1, localMem[982], 2);
              ip = 2245;
      end

       2245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1004] = heapMem[localMem[981]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2246;
      end

       2246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1005] = heapMem[localMem[981]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2247;
      end

       2247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1006] = heapMem[localMem[1005]*6 + localMem[1004]];
              updateArrayLength(2, 0, 0);
              ip = 2248;
      end

       2248 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1006] != localMem[974] ? 2267 : 2249;
      end

       2249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1007] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2250;
      end

       2250 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1008] = heapMem[localMem[1007]*6 + localMem[979]];
              updateArrayLength(2, 0, 0);
              ip = 2251;
      end

       2251 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1009] = heapMem[localMem[981]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2252;
      end

       2252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1009]*6 + localMem[1004]] = localMem[1008];
              updateArrayLength(1, localMem[1009], localMem[1004]);
              ip = 2253;
      end

       2253 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1010] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2254;
      end

       2254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1011] = heapMem[localMem[1010]*6 + localMem[979]];
              updateArrayLength(2, 0, 0);
              ip = 2255;
      end

       2255 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1012] = heapMem[localMem[981]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2256;
      end

       2256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1012]*6 + localMem[1004]] = localMem[1011];
              updateArrayLength(1, localMem[1012], localMem[1004]);
              ip = 2257;
      end

       2257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1013] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2258;
      end

       2258 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1013]] = localMem[979];
              ip = 2259;
      end

       2259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1014] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2260;
      end

       2260 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1014]] = localMem[979];
              ip = 2261;
      end

       2261 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1015] = localMem[1004] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2262;
      end

       2262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[981]*6 + 0] = localMem[1015];
              updateArrayLength(1, localMem[981], 0);
              ip = 2263;
      end

       2263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1016] = heapMem[localMem[981]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2264;
      end

       2264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1016]*6 + localMem[1015]] = localMem[982];
              updateArrayLength(1, localMem[1016], localMem[1015]);
              ip = 2265;
      end

       2265 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2405;
      end

       2266 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2289;
      end

       2267 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2268;
      end

       2268 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 2269;
      end

       2269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1017] = heapMem[localMem[981]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2270;
      end

       2270 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1018] = 0; k = arraySizes[localMem[1017]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1017] * NArea + i] == localMem[974]) localMem[1018] = i + 1;
              end
              ip = 2271;
      end

       2271 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1018] = localMem[1018] - 1;
              updateArrayLength(2, 0, 0);
              ip = 2272;
      end

       2272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1019] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2273;
      end

       2273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1020] = heapMem[localMem[1019]*6 + localMem[979]];
              updateArrayLength(2, 0, 0);
              ip = 2274;
      end

       2274 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1021] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2275;
      end

       2275 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1022] = heapMem[localMem[1021]*6 + localMem[979]];
              updateArrayLength(2, 0, 0);
              ip = 2276;
      end

       2276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1023] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2277;
      end

       2277 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1023]] = localMem[979];
              ip = 2278;
      end

       2278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1024] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2279;
      end

       2279 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1024]] = localMem[979];
              ip = 2280;
      end

       2280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1025] = heapMem[localMem[981]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2281;
      end

       2281 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1025] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1018], localMem[1025], arraySizes[localMem[1025]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1018] && i <= arraySizes[localMem[1025]]) begin
                  heapMem[NArea * localMem[1025] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1025] + localMem[1018]] = localMem[1020];                                    // Insert new value
              arraySizes[localMem[1025]] = arraySizes[localMem[1025]] + 1;                              // Increase array size
              ip = 2282;
      end

       2282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1026] = heapMem[localMem[981]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2283;
      end

       2283 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1026] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1018], localMem[1026], arraySizes[localMem[1026]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1018] && i <= arraySizes[localMem[1026]]) begin
                  heapMem[NArea * localMem[1026] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1026] + localMem[1018]] = localMem[1022];                                    // Insert new value
              arraySizes[localMem[1026]] = arraySizes[localMem[1026]] + 1;                              // Increase array size
              ip = 2284;
      end

       2284 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1027] = heapMem[localMem[981]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2285;
      end

       2285 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1028] = localMem[1018] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2286;
      end

       2286 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1027] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1028], localMem[1027], arraySizes[localMem[1027]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1028] && i <= arraySizes[localMem[1027]]) begin
                  heapMem[NArea * localMem[1027] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1027] + localMem[1028]] = localMem[982];                                    // Insert new value
              arraySizes[localMem[1027]] = arraySizes[localMem[1027]] + 1;                              // Increase array size
              ip = 2287;
      end

       2287 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[981]*6 + 0] = heapMem[localMem[981]*6 + 0] + 1;
              updateArrayLength(1, localMem[981], 0);
              ip = 2288;
      end

       2288 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2405;
      end

       2289 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2290;
      end

       2290 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2291;
      end

       2291 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1029] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1029] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1029]] = 0;
              ip = 2292;
      end

       2292 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 0] = localMem[979];
              updateArrayLength(1, localMem[1029], 0);
              ip = 2293;
      end

       2293 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 2] = 0;
              updateArrayLength(1, localMem[1029], 2);
              ip = 2294;
      end

       2294 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1030] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1030] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1030]] = 0;
              ip = 2295;
      end

       2295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 4] = localMem[1030];
              updateArrayLength(1, localMem[1029], 4);
              ip = 2296;
      end

       2296 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1031] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1031] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1031]] = 0;
              ip = 2297;
      end

       2297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 5] = localMem[1031];
              updateArrayLength(1, localMem[1029], 5);
              ip = 2298;
      end

       2298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 6] = 0;
              updateArrayLength(1, localMem[1029], 6);
              ip = 2299;
      end

       2299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 3] = localMem[977];
              updateArrayLength(1, localMem[1029], 3);
              ip = 2300;
      end

       2300 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[977]*6 + 1] = heapMem[localMem[977]*6 + 1] + 1;
              updateArrayLength(1, localMem[977], 1);
              ip = 2301;
      end

       2301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 1] = heapMem[localMem[977]*6 + 1];
              updateArrayLength(1, localMem[1029], 1);
              ip = 2302;
      end

       2302 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1032] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1032] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1032]] = 0;
              ip = 2303;
      end

       2303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 0] = localMem[979];
              updateArrayLength(1, localMem[1032], 0);
              ip = 2304;
      end

       2304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 2] = 0;
              updateArrayLength(1, localMem[1032], 2);
              ip = 2305;
      end

       2305 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1033] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1033] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1033]] = 0;
              ip = 2306;
      end

       2306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 4] = localMem[1033];
              updateArrayLength(1, localMem[1032], 4);
              ip = 2307;
      end

       2307 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1034] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1034] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1034]] = 0;
              ip = 2308;
      end

       2308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 5] = localMem[1034];
              updateArrayLength(1, localMem[1032], 5);
              ip = 2309;
      end

       2309 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 6] = 0;
              updateArrayLength(1, localMem[1032], 6);
              ip = 2310;
      end

       2310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 3] = localMem[977];
              updateArrayLength(1, localMem[1032], 3);
              ip = 2311;
      end

       2311 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[977]*6 + 1] = heapMem[localMem[977]*6 + 1] + 1;
              updateArrayLength(1, localMem[977], 1);
              ip = 2312;
      end

       2312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 1] = heapMem[localMem[977]*6 + 1];
              updateArrayLength(1, localMem[1032], 1);
              ip = 2313;
      end

       2313 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1035] = !heapMem[localMem[974]*6 + 6];
              ip = 2314;
      end

       2314 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1035] != 0 ? 2366 : 2315;
      end

       2315 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1036] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1036] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1036]] = 0;
              ip = 2316;
      end

       2316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 6] = localMem[1036];
              updateArrayLength(1, localMem[1029], 6);
              ip = 2317;
      end

       2317 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1037] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1037] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1037]] = 0;
              ip = 2318;
      end

       2318 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 6] = localMem[1037];
              updateArrayLength(1, localMem[1032], 6);
              ip = 2319;
      end

       2319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1038] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2320;
      end

       2320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1039] = heapMem[localMem[1029]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2321;
      end

       2321 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1039] + 0 + i] = heapMem[NArea * localMem[1038] + 0 + i];
                  updateArrayLength(1, localMem[1039], 0 + i);
                end
              end
              ip = 2322;
      end

       2322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1040] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2323;
      end

       2323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1041] = heapMem[localMem[1029]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2324;
      end

       2324 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1041] + 0 + i] = heapMem[NArea * localMem[1040] + 0 + i];
                  updateArrayLength(1, localMem[1041], 0 + i);
                end
              end
              ip = 2325;
      end

       2325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1042] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2326;
      end

       2326 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1043] = heapMem[localMem[1029]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2327;
      end

       2327 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1044] = localMem[979] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2328;
      end

       2328 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1044]) begin
                  heapMem[NArea * localMem[1043] + 0 + i] = heapMem[NArea * localMem[1042] + 0 + i];
                  updateArrayLength(1, localMem[1043], 0 + i);
                end
              end
              ip = 2329;
      end

       2329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1045] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2330;
      end

       2330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1046] = heapMem[localMem[1032]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2331;
      end

       2331 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1046] + 0 + i] = heapMem[NArea * localMem[1045] + localMem[980] + i];
                  updateArrayLength(1, localMem[1046], 0 + i);
                end
              end
              ip = 2332;
      end

       2332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1047] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2333;
      end

       2333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1048] = heapMem[localMem[1032]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2334;
      end

       2334 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1048] + 0 + i] = heapMem[NArea * localMem[1047] + localMem[980] + i];
                  updateArrayLength(1, localMem[1048], 0 + i);
                end
              end
              ip = 2335;
      end

       2335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1049] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2336;
      end

       2336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1050] = heapMem[localMem[1032]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2337;
      end

       2337 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1051] = localMem[979] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2338;
      end

       2338 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1051]) begin
                  heapMem[NArea * localMem[1050] + 0 + i] = heapMem[NArea * localMem[1049] + localMem[980] + i];
                  updateArrayLength(1, localMem[1050], 0 + i);
                end
              end
              ip = 2339;
      end

       2339 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1052] = heapMem[localMem[1029]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2340;
      end

       2340 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1053] = localMem[1052] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2341;
      end

       2341 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1054] = heapMem[localMem[1029]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2342;
      end

       2342 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2343;
      end

       2343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1055] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2344;
      end

       2344 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2345;
      end

       2345 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1055] >= localMem[1053] ? 2351 : 2346;
      end

       2346 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1056] = heapMem[localMem[1054]*6 + localMem[1055]];
              updateArrayLength(2, 0, 0);
              ip = 2347;
      end

       2347 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1056]*6 + 2] = localMem[1029];
              updateArrayLength(1, localMem[1056], 2);
              ip = 2348;
      end

       2348 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2349;
      end

       2349 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1055] = localMem[1055] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2350;
      end

       2350 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2344;
      end

       2351 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2352;
      end

       2352 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1057] = heapMem[localMem[1032]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2353;
      end

       2353 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1058] = localMem[1057] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2354;
      end

       2354 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1059] = heapMem[localMem[1032]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2355;
      end

       2355 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2356;
      end

       2356 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1060] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2357;
      end

       2357 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2358;
      end

       2358 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1060] >= localMem[1058] ? 2364 : 2359;
      end

       2359 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1061] = heapMem[localMem[1059]*6 + localMem[1060]];
              updateArrayLength(2, 0, 0);
              ip = 2360;
      end

       2360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1061]*6 + 2] = localMem[1032];
              updateArrayLength(1, localMem[1061], 2);
              ip = 2361;
      end

       2361 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2362;
      end

       2362 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1060] = localMem[1060] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2363;
      end

       2363 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2357;
      end

       2364 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2365;
      end

       2365 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2381;
      end

       2366 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2367;
      end

       2367 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1062] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1062] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1062]] = 0;
              ip = 2368;
      end

       2368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[974]*6 + 6] = localMem[1062];
              updateArrayLength(1, localMem[974], 6);
              ip = 2369;
      end

       2369 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1063] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2370;
      end

       2370 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1064] = heapMem[localMem[1029]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2371;
      end

       2371 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1064] + 0 + i] = heapMem[NArea * localMem[1063] + 0 + i];
                  updateArrayLength(1, localMem[1064], 0 + i);
                end
              end
              ip = 2372;
      end

       2372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1065] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2373;
      end

       2373 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1066] = heapMem[localMem[1029]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2374;
      end

       2374 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1066] + 0 + i] = heapMem[NArea * localMem[1065] + 0 + i];
                  updateArrayLength(1, localMem[1066], 0 + i);
                end
              end
              ip = 2375;
      end

       2375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1067] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2376;
      end

       2376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1068] = heapMem[localMem[1032]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2377;
      end

       2377 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1068] + 0 + i] = heapMem[NArea * localMem[1067] + localMem[980] + i];
                  updateArrayLength(1, localMem[1068], 0 + i);
                end
              end
              ip = 2378;
      end

       2378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1069] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2379;
      end

       2379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1070] = heapMem[localMem[1032]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2380;
      end

       2380 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[979]) begin
                  heapMem[NArea * localMem[1070] + 0 + i] = heapMem[NArea * localMem[1069] + localMem[980] + i];
                  updateArrayLength(1, localMem[1070], 0 + i);
                end
              end
              ip = 2381;
      end

       2381 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2382;
      end

       2382 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1029]*6 + 2] = localMem[974];
              updateArrayLength(1, localMem[1029], 2);
              ip = 2383;
      end

       2383 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1032]*6 + 2] = localMem[974];
              updateArrayLength(1, localMem[1032], 2);
              ip = 2384;
      end

       2384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1071] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2385;
      end

       2385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1072] = heapMem[localMem[1071]*6 + localMem[979]];
              updateArrayLength(2, 0, 0);
              ip = 2386;
      end

       2386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1073] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2387;
      end

       2387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1074] = heapMem[localMem[1073]*6 + localMem[979]];
              updateArrayLength(2, 0, 0);
              ip = 2388;
      end

       2388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1075] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2389;
      end

       2389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1075]*6 + 0] = localMem[1072];
              updateArrayLength(1, localMem[1075], 0);
              ip = 2390;
      end

       2390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1076] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2391;
      end

       2391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1076]*6 + 0] = localMem[1074];
              updateArrayLength(1, localMem[1076], 0);
              ip = 2392;
      end

       2392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1077] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2393;
      end

       2393 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1077]*6 + 0] = localMem[1029];
              updateArrayLength(1, localMem[1077], 0);
              ip = 2394;
      end

       2394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1078] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2395;
      end

       2395 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1078]*6 + 1] = localMem[1032];
              updateArrayLength(1, localMem[1078], 1);
              ip = 2396;
      end

       2396 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[974]*6 + 0] = 1;
              updateArrayLength(1, localMem[974], 0);
              ip = 2397;
      end

       2397 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1079] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2398;
      end

       2398 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1079]] = 1;
              ip = 2399;
      end

       2399 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1080] = heapMem[localMem[974]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2400;
      end

       2400 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1080]] = 1;
              ip = 2401;
      end

       2401 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1081] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2402;
      end

       2402 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1081]] = 2;
              ip = 2403;
      end

       2403 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2405;
      end

       2404 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2410;
      end

       2405 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2406;
      end

       2406 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[975] = 1;
              updateArrayLength(2, 0, 0);
              ip = 2407;
      end

       2407 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2410;
      end

       2408 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2409;
      end

       2409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[975] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2410;
      end

       2410 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2411;
      end

       2411 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2412;
      end

       2412 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2413;
      end

       2413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1082] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2414;
      end

       2414 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2415;
      end

       2415 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1082] >= 99 ? 2913 : 2416;
      end

       2416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1083] = heapMem[localMem[974]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2417;
      end

       2417 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1084] = localMem[1083] - 1;
              updateArrayLength(2, 0, 0);
              ip = 2418;
      end

       2418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1085] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2419;
      end

       2419 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1086] = heapMem[localMem[1085]*6 + localMem[1084]];
              updateArrayLength(2, 0, 0);
              ip = 2420;
      end

       2420 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 3 <= localMem[1086] ? 2661 : 2421;
      end

       2421 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1087] = !heapMem[localMem[974]*6 + 6];
              ip = 2422;
      end

       2422 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1087] == 0 ? 2427 : 2423;
      end

       2423 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 0] = localMem[974];
              updateArrayLength(1, localMem[951], 0);
              ip = 2424;
      end

       2424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 1] = 2;
              updateArrayLength(1, localMem[951], 1);
              ip = 2425;
      end

       2425 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[951]*6 + 2] = localMem[1083] - 1;
              updateArrayLength(1, localMem[951], 2);
              ip = 2426;
      end

       2426 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2917;
      end

       2427 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2428;
      end

       2428 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1088] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2429;
      end

       2429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1089] = heapMem[localMem[1088]*6 + localMem[1083]];
              updateArrayLength(2, 0, 0);
              ip = 2430;
      end

       2430 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2431;
      end

       2431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1091] = heapMem[localMem[1089]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2432;
      end

       2432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1092] = heapMem[localMem[1089]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2433;
      end

       2433 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1093] = heapMem[localMem[1092]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2434;
      end

       2434 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1091] <  localMem[1093] ? 2654 : 2435;
      end

       2435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1094] = localMem[1093];
              updateArrayLength(2, 0, 0);
              ip = 2436;
      end

       2436 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1094] = localMem[1094] >> 1;
              ip = 2437;
      end

       2437 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1095] = localMem[1094] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2438;
      end

       2438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1096] = heapMem[localMem[1089]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2439;
      end

       2439 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1096] == 0 ? 2536 : 2440;
      end

       2440 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1097] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1097] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1097]] = 0;
              ip = 2441;
      end

       2441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 0] = localMem[1094];
              updateArrayLength(1, localMem[1097], 0);
              ip = 2442;
      end

       2442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 2] = 0;
              updateArrayLength(1, localMem[1097], 2);
              ip = 2443;
      end

       2443 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1098] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1098] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1098]] = 0;
              ip = 2444;
      end

       2444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 4] = localMem[1098];
              updateArrayLength(1, localMem[1097], 4);
              ip = 2445;
      end

       2445 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1099] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1099] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1099]] = 0;
              ip = 2446;
      end

       2446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 5] = localMem[1099];
              updateArrayLength(1, localMem[1097], 5);
              ip = 2447;
      end

       2447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 6] = 0;
              updateArrayLength(1, localMem[1097], 6);
              ip = 2448;
      end

       2448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 3] = localMem[1092];
              updateArrayLength(1, localMem[1097], 3);
              ip = 2449;
      end

       2449 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1092]*6 + 1] = heapMem[localMem[1092]*6 + 1] + 1;
              updateArrayLength(1, localMem[1092], 1);
              ip = 2450;
      end

       2450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 1] = heapMem[localMem[1092]*6 + 1];
              updateArrayLength(1, localMem[1097], 1);
              ip = 2451;
      end

       2451 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1100] = !heapMem[localMem[1089]*6 + 6];
              ip = 2452;
      end

       2452 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1100] != 0 ? 2481 : 2453;
      end

       2453 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1101] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1101] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1101]] = 0;
              ip = 2454;
      end

       2454 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 6] = localMem[1101];
              updateArrayLength(1, localMem[1097], 6);
              ip = 2455;
      end

       2455 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1102] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2456;
      end

       2456 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1103] = heapMem[localMem[1097]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2457;
      end

       2457 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1103] + 0 + i] = heapMem[NArea * localMem[1102] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1103], 0 + i);
                end
              end
              ip = 2458;
      end

       2458 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1104] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2459;
      end

       2459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1105] = heapMem[localMem[1097]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2460;
      end

       2460 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1105] + 0 + i] = heapMem[NArea * localMem[1104] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1105], 0 + i);
                end
              end
              ip = 2461;
      end

       2461 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1106] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2462;
      end

       2462 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1107] = heapMem[localMem[1097]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2463;
      end

       2463 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1108] = localMem[1094] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2464;
      end

       2464 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1108]) begin
                  heapMem[NArea * localMem[1107] + 0 + i] = heapMem[NArea * localMem[1106] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1107], 0 + i);
                end
              end
              ip = 2465;
      end

       2465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1109] = heapMem[localMem[1097]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2466;
      end

       2466 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1110] = localMem[1109] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2467;
      end

       2467 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1111] = heapMem[localMem[1097]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2468;
      end

       2468 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2469;
      end

       2469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1112] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2470;
      end

       2470 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2471;
      end

       2471 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1112] >= localMem[1110] ? 2477 : 2472;
      end

       2472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1113] = heapMem[localMem[1111]*6 + localMem[1112]];
              updateArrayLength(2, 0, 0);
              ip = 2473;
      end

       2473 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1113]*6 + 2] = localMem[1097];
              updateArrayLength(1, localMem[1113], 2);
              ip = 2474;
      end

       2474 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2475;
      end

       2475 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1112] = localMem[1112] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2476;
      end

       2476 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2470;
      end

       2477 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2478;
      end

       2478 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1114] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2479;
      end

       2479 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1114]] = localMem[1095];
              ip = 2480;
      end

       2480 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2488;
      end

       2481 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2482;
      end

       2482 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1115] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2483;
      end

       2483 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1116] = heapMem[localMem[1097]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2484;
      end

       2484 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1116] + 0 + i] = heapMem[NArea * localMem[1115] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1116], 0 + i);
                end
              end
              ip = 2485;
      end

       2485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1117] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2486;
      end

       2486 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1118] = heapMem[localMem[1097]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2487;
      end

       2487 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1118] + 0 + i] = heapMem[NArea * localMem[1117] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1118], 0 + i);
                end
              end
              ip = 2488;
      end

       2488 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2489;
      end

       2489 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1089]*6 + 0] = localMem[1094];
              updateArrayLength(1, localMem[1089], 0);
              ip = 2490;
      end

       2490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1097]*6 + 2] = localMem[1096];
              updateArrayLength(1, localMem[1097], 2);
              ip = 2491;
      end

       2491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1119] = heapMem[localMem[1096]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2492;
      end

       2492 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1120] = heapMem[localMem[1096]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2493;
      end

       2493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1121] = heapMem[localMem[1120]*6 + localMem[1119]];
              updateArrayLength(2, 0, 0);
              ip = 2494;
      end

       2494 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1121] != localMem[1089] ? 2513 : 2495;
      end

       2495 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1122] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2496;
      end

       2496 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1123] = heapMem[localMem[1122]*6 + localMem[1094]];
              updateArrayLength(2, 0, 0);
              ip = 2497;
      end

       2497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1124] = heapMem[localMem[1096]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2498;
      end

       2498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1124]*6 + localMem[1119]] = localMem[1123];
              updateArrayLength(1, localMem[1124], localMem[1119]);
              ip = 2499;
      end

       2499 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1125] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2500;
      end

       2500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1126] = heapMem[localMem[1125]*6 + localMem[1094]];
              updateArrayLength(2, 0, 0);
              ip = 2501;
      end

       2501 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1127] = heapMem[localMem[1096]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2502;
      end

       2502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1127]*6 + localMem[1119]] = localMem[1126];
              updateArrayLength(1, localMem[1127], localMem[1119]);
              ip = 2503;
      end

       2503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1128] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2504;
      end

       2504 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1128]] = localMem[1094];
              ip = 2505;
      end

       2505 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1129] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2506;
      end

       2506 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1129]] = localMem[1094];
              ip = 2507;
      end

       2507 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1130] = localMem[1119] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2508;
      end

       2508 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1096]*6 + 0] = localMem[1130];
              updateArrayLength(1, localMem[1096], 0);
              ip = 2509;
      end

       2509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1131] = heapMem[localMem[1096]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2510;
      end

       2510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1131]*6 + localMem[1130]] = localMem[1097];
              updateArrayLength(1, localMem[1131], localMem[1130]);
              ip = 2511;
      end

       2511 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2651;
      end

       2512 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2535;
      end

       2513 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2514;
      end

       2514 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 2515;
      end

       2515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1132] = heapMem[localMem[1096]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2516;
      end

       2516 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1133] = 0; k = arraySizes[localMem[1132]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1132] * NArea + i] == localMem[1089]) localMem[1133] = i + 1;
              end
              ip = 2517;
      end

       2517 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1133] = localMem[1133] - 1;
              updateArrayLength(2, 0, 0);
              ip = 2518;
      end

       2518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1134] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2519;
      end

       2519 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1135] = heapMem[localMem[1134]*6 + localMem[1094]];
              updateArrayLength(2, 0, 0);
              ip = 2520;
      end

       2520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1136] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2521;
      end

       2521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1137] = heapMem[localMem[1136]*6 + localMem[1094]];
              updateArrayLength(2, 0, 0);
              ip = 2522;
      end

       2522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1138] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2523;
      end

       2523 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1138]] = localMem[1094];
              ip = 2524;
      end

       2524 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1139] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2525;
      end

       2525 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1139]] = localMem[1094];
              ip = 2526;
      end

       2526 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1140] = heapMem[localMem[1096]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2527;
      end

       2527 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1140] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1133], localMem[1140], arraySizes[localMem[1140]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1133] && i <= arraySizes[localMem[1140]]) begin
                  heapMem[NArea * localMem[1140] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1140] + localMem[1133]] = localMem[1135];                                    // Insert new value
              arraySizes[localMem[1140]] = arraySizes[localMem[1140]] + 1;                              // Increase array size
              ip = 2528;
      end

       2528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1141] = heapMem[localMem[1096]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2529;
      end

       2529 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1141] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1133], localMem[1141], arraySizes[localMem[1141]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1133] && i <= arraySizes[localMem[1141]]) begin
                  heapMem[NArea * localMem[1141] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1141] + localMem[1133]] = localMem[1137];                                    // Insert new value
              arraySizes[localMem[1141]] = arraySizes[localMem[1141]] + 1;                              // Increase array size
              ip = 2530;
      end

       2530 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1142] = heapMem[localMem[1096]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2531;
      end

       2531 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1143] = localMem[1133] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2532;
      end

       2532 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1142] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1143], localMem[1142], arraySizes[localMem[1142]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1143] && i <= arraySizes[localMem[1142]]) begin
                  heapMem[NArea * localMem[1142] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1142] + localMem[1143]] = localMem[1097];                                    // Insert new value
              arraySizes[localMem[1142]] = arraySizes[localMem[1142]] + 1;                              // Increase array size
              ip = 2533;
      end

       2533 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1096]*6 + 0] = heapMem[localMem[1096]*6 + 0] + 1;
              updateArrayLength(1, localMem[1096], 0);
              ip = 2534;
      end

       2534 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2651;
      end

       2535 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2536;
      end

       2536 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2537;
      end

       2537 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1144] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1144] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1144]] = 0;
              ip = 2538;
      end

       2538 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 0] = localMem[1094];
              updateArrayLength(1, localMem[1144], 0);
              ip = 2539;
      end

       2539 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 2] = 0;
              updateArrayLength(1, localMem[1144], 2);
              ip = 2540;
      end

       2540 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1145] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1145] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1145]] = 0;
              ip = 2541;
      end

       2541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 4] = localMem[1145];
              updateArrayLength(1, localMem[1144], 4);
              ip = 2542;
      end

       2542 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1146] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1146] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1146]] = 0;
              ip = 2543;
      end

       2543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 5] = localMem[1146];
              updateArrayLength(1, localMem[1144], 5);
              ip = 2544;
      end

       2544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 6] = 0;
              updateArrayLength(1, localMem[1144], 6);
              ip = 2545;
      end

       2545 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 3] = localMem[1092];
              updateArrayLength(1, localMem[1144], 3);
              ip = 2546;
      end

       2546 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1092]*6 + 1] = heapMem[localMem[1092]*6 + 1] + 1;
              updateArrayLength(1, localMem[1092], 1);
              ip = 2547;
      end

       2547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 1] = heapMem[localMem[1092]*6 + 1];
              updateArrayLength(1, localMem[1144], 1);
              ip = 2548;
      end

       2548 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1147] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1147] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1147]] = 0;
              ip = 2549;
      end

       2549 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 0] = localMem[1094];
              updateArrayLength(1, localMem[1147], 0);
              ip = 2550;
      end

       2550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 2] = 0;
              updateArrayLength(1, localMem[1147], 2);
              ip = 2551;
      end

       2551 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1148] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1148] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1148]] = 0;
              ip = 2552;
      end

       2552 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 4] = localMem[1148];
              updateArrayLength(1, localMem[1147], 4);
              ip = 2553;
      end

       2553 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1149] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1149] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1149]] = 0;
              ip = 2554;
      end

       2554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 5] = localMem[1149];
              updateArrayLength(1, localMem[1147], 5);
              ip = 2555;
      end

       2555 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 6] = 0;
              updateArrayLength(1, localMem[1147], 6);
              ip = 2556;
      end

       2556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 3] = localMem[1092];
              updateArrayLength(1, localMem[1147], 3);
              ip = 2557;
      end

       2557 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1092]*6 + 1] = heapMem[localMem[1092]*6 + 1] + 1;
              updateArrayLength(1, localMem[1092], 1);
              ip = 2558;
      end

       2558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 1] = heapMem[localMem[1092]*6 + 1];
              updateArrayLength(1, localMem[1147], 1);
              ip = 2559;
      end

       2559 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1150] = !heapMem[localMem[1089]*6 + 6];
              ip = 2560;
      end

       2560 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1150] != 0 ? 2612 : 2561;
      end

       2561 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1151] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1151] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1151]] = 0;
              ip = 2562;
      end

       2562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 6] = localMem[1151];
              updateArrayLength(1, localMem[1144], 6);
              ip = 2563;
      end

       2563 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1152] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1152] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1152]] = 0;
              ip = 2564;
      end

       2564 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 6] = localMem[1152];
              updateArrayLength(1, localMem[1147], 6);
              ip = 2565;
      end

       2565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1153] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2566;
      end

       2566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1154] = heapMem[localMem[1144]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2567;
      end

       2567 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1154] + 0 + i] = heapMem[NArea * localMem[1153] + 0 + i];
                  updateArrayLength(1, localMem[1154], 0 + i);
                end
              end
              ip = 2568;
      end

       2568 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1155] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2569;
      end

       2569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1156] = heapMem[localMem[1144]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2570;
      end

       2570 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1156] + 0 + i] = heapMem[NArea * localMem[1155] + 0 + i];
                  updateArrayLength(1, localMem[1156], 0 + i);
                end
              end
              ip = 2571;
      end

       2571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1157] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2572;
      end

       2572 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1158] = heapMem[localMem[1144]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2573;
      end

       2573 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1159] = localMem[1094] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2574;
      end

       2574 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1159]) begin
                  heapMem[NArea * localMem[1158] + 0 + i] = heapMem[NArea * localMem[1157] + 0 + i];
                  updateArrayLength(1, localMem[1158], 0 + i);
                end
              end
              ip = 2575;
      end

       2575 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1160] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2576;
      end

       2576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1161] = heapMem[localMem[1147]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2577;
      end

       2577 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1161] + 0 + i] = heapMem[NArea * localMem[1160] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1161], 0 + i);
                end
              end
              ip = 2578;
      end

       2578 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1162] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2579;
      end

       2579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1163] = heapMem[localMem[1147]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2580;
      end

       2580 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1163] + 0 + i] = heapMem[NArea * localMem[1162] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1163], 0 + i);
                end
              end
              ip = 2581;
      end

       2581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1164] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2582;
      end

       2582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1165] = heapMem[localMem[1147]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2583;
      end

       2583 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1166] = localMem[1094] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2584;
      end

       2584 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1166]) begin
                  heapMem[NArea * localMem[1165] + 0 + i] = heapMem[NArea * localMem[1164] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1165], 0 + i);
                end
              end
              ip = 2585;
      end

       2585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1167] = heapMem[localMem[1144]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2586;
      end

       2586 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1168] = localMem[1167] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2587;
      end

       2587 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1169] = heapMem[localMem[1144]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2588;
      end

       2588 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2589;
      end

       2589 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1170] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2590;
      end

       2590 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2591;
      end

       2591 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1170] >= localMem[1168] ? 2597 : 2592;
      end

       2592 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1171] = heapMem[localMem[1169]*6 + localMem[1170]];
              updateArrayLength(2, 0, 0);
              ip = 2593;
      end

       2593 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1171]*6 + 2] = localMem[1144];
              updateArrayLength(1, localMem[1171], 2);
              ip = 2594;
      end

       2594 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2595;
      end

       2595 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1170] = localMem[1170] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2596;
      end

       2596 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2590;
      end

       2597 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2598;
      end

       2598 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1172] = heapMem[localMem[1147]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2599;
      end

       2599 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1173] = localMem[1172] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2600;
      end

       2600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1174] = heapMem[localMem[1147]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2601;
      end

       2601 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2602;
      end

       2602 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1175] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2603;
      end

       2603 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2604;
      end

       2604 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1175] >= localMem[1173] ? 2610 : 2605;
      end

       2605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1176] = heapMem[localMem[1174]*6 + localMem[1175]];
              updateArrayLength(2, 0, 0);
              ip = 2606;
      end

       2606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1176]*6 + 2] = localMem[1147];
              updateArrayLength(1, localMem[1176], 2);
              ip = 2607;
      end

       2607 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2608;
      end

       2608 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1175] = localMem[1175] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2609;
      end

       2609 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2603;
      end

       2610 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2611;
      end

       2611 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2627;
      end

       2612 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2613;
      end

       2613 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1177] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1177] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1177]] = 0;
              ip = 2614;
      end

       2614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1089]*6 + 6] = localMem[1177];
              updateArrayLength(1, localMem[1089], 6);
              ip = 2615;
      end

       2615 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1178] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2616;
      end

       2616 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1179] = heapMem[localMem[1144]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2617;
      end

       2617 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1179] + 0 + i] = heapMem[NArea * localMem[1178] + 0 + i];
                  updateArrayLength(1, localMem[1179], 0 + i);
                end
              end
              ip = 2618;
      end

       2618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1180] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2619;
      end

       2619 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1181] = heapMem[localMem[1144]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2620;
      end

       2620 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1181] + 0 + i] = heapMem[NArea * localMem[1180] + 0 + i];
                  updateArrayLength(1, localMem[1181], 0 + i);
                end
              end
              ip = 2621;
      end

       2621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1182] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2622;
      end

       2622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1183] = heapMem[localMem[1147]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2623;
      end

       2623 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1183] + 0 + i] = heapMem[NArea * localMem[1182] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1183], 0 + i);
                end
              end
              ip = 2624;
      end

       2624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1184] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2625;
      end

       2625 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1185] = heapMem[localMem[1147]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2626;
      end

       2626 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1094]) begin
                  heapMem[NArea * localMem[1185] + 0 + i] = heapMem[NArea * localMem[1184] + localMem[1095] + i];
                  updateArrayLength(1, localMem[1185], 0 + i);
                end
              end
              ip = 2627;
      end

       2627 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2628;
      end

       2628 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1144]*6 + 2] = localMem[1089];
              updateArrayLength(1, localMem[1144], 2);
              ip = 2629;
      end

       2629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1147]*6 + 2] = localMem[1089];
              updateArrayLength(1, localMem[1147], 2);
              ip = 2630;
      end

       2630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1186] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2631;
      end

       2631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1187] = heapMem[localMem[1186]*6 + localMem[1094]];
              updateArrayLength(2, 0, 0);
              ip = 2632;
      end

       2632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1188] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2633;
      end

       2633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1189] = heapMem[localMem[1188]*6 + localMem[1094]];
              updateArrayLength(2, 0, 0);
              ip = 2634;
      end

       2634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1190] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2635;
      end

       2635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1190]*6 + 0] = localMem[1187];
              updateArrayLength(1, localMem[1190], 0);
              ip = 2636;
      end

       2636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1191] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2637;
      end

       2637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1191]*6 + 0] = localMem[1189];
              updateArrayLength(1, localMem[1191], 0);
              ip = 2638;
      end

       2638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1192] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2639;
      end

       2639 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1192]*6 + 0] = localMem[1144];
              updateArrayLength(1, localMem[1192], 0);
              ip = 2640;
      end

       2640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1193] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2641;
      end

       2641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1193]*6 + 1] = localMem[1147];
              updateArrayLength(1, localMem[1193], 1);
              ip = 2642;
      end

       2642 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1089]*6 + 0] = 1;
              updateArrayLength(1, localMem[1089], 0);
              ip = 2643;
      end

       2643 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1194] = heapMem[localMem[1089]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2644;
      end

       2644 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1194]] = 1;
              ip = 2645;
      end

       2645 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1195] = heapMem[localMem[1089]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2646;
      end

       2646 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1195]] = 1;
              ip = 2647;
      end

       2647 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1196] = heapMem[localMem[1089]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2648;
      end

       2648 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1196]] = 2;
              ip = 2649;
      end

       2649 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2651;
      end

       2650 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2656;
      end

       2651 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2652;
      end

       2652 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1090] = 1;
              updateArrayLength(2, 0, 0);
              ip = 2653;
      end

       2653 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2656;
      end

       2654 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2655;
      end

       2655 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1090] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2656;
      end

       2656 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2657;
      end

       2657 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1090] != 0 ? 2659 : 2658;
      end

       2658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[974] = localMem[1089];
              updateArrayLength(2, 0, 0);
              ip = 2659;
      end

       2659 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2660;
      end

       2660 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2910;
      end

       2661 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2662;
      end

       2662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1197] = heapMem[localMem[974]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2663;
      end

       2663 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1198] = 0; k = arraySizes[localMem[1197]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1197] * NArea + i] == 3) localMem[1198] = i + 1;
              end
              ip = 2664;
      end

       2664 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1198] == 0 ? 2669 : 2665;
      end

       2665 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 0] = localMem[974];
              updateArrayLength(1, localMem[951], 0);
              ip = 2666;
      end

       2666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 1] = 1;
              updateArrayLength(1, localMem[951], 1);
              ip = 2667;
      end

       2667 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[951]*6 + 2] = localMem[1198] - 1;
              updateArrayLength(1, localMem[951], 2);
              ip = 2668;
      end

       2668 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2917;
      end

       2669 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2670;
      end

       2670 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[1197]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1197] * NArea + i] < 3) j = j + 1;
              end
              localMem[1199] = j;
              ip = 2671;
      end

       2671 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1200] = !heapMem[localMem[974]*6 + 6];
              ip = 2672;
      end

       2672 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1200] == 0 ? 2677 : 2673;
      end

       2673 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 0] = localMem[974];
              updateArrayLength(1, localMem[951], 0);
              ip = 2674;
      end

       2674 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 1] = 0;
              updateArrayLength(1, localMem[951], 1);
              ip = 2675;
      end

       2675 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[951]*6 + 2] = localMem[1199];
              updateArrayLength(1, localMem[951], 2);
              ip = 2676;
      end

       2676 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2917;
      end

       2677 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2678;
      end

       2678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1201] = heapMem[localMem[974]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2679;
      end

       2679 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1202] = heapMem[localMem[1201]*6 + localMem[1199]];
              updateArrayLength(2, 0, 0);
              ip = 2680;
      end

       2680 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2681;
      end

       2681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1204] = heapMem[localMem[1202]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2682;
      end

       2682 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1205] = heapMem[localMem[1202]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2683;
      end

       2683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1206] = heapMem[localMem[1205]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2684;
      end

       2684 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1204] <  localMem[1206] ? 2904 : 2685;
      end

       2685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1207] = localMem[1206];
              updateArrayLength(2, 0, 0);
              ip = 2686;
      end

       2686 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1207] = localMem[1207] >> 1;
              ip = 2687;
      end

       2687 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1208] = localMem[1207] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2688;
      end

       2688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1209] = heapMem[localMem[1202]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2689;
      end

       2689 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1209] == 0 ? 2786 : 2690;
      end

       2690 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1210] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1210] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1210]] = 0;
              ip = 2691;
      end

       2691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 0] = localMem[1207];
              updateArrayLength(1, localMem[1210], 0);
              ip = 2692;
      end

       2692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 2] = 0;
              updateArrayLength(1, localMem[1210], 2);
              ip = 2693;
      end

       2693 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1211] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1211] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1211]] = 0;
              ip = 2694;
      end

       2694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 4] = localMem[1211];
              updateArrayLength(1, localMem[1210], 4);
              ip = 2695;
      end

       2695 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1212] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1212] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1212]] = 0;
              ip = 2696;
      end

       2696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 5] = localMem[1212];
              updateArrayLength(1, localMem[1210], 5);
              ip = 2697;
      end

       2697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 6] = 0;
              updateArrayLength(1, localMem[1210], 6);
              ip = 2698;
      end

       2698 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 3] = localMem[1205];
              updateArrayLength(1, localMem[1210], 3);
              ip = 2699;
      end

       2699 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1205]*6 + 1] = heapMem[localMem[1205]*6 + 1] + 1;
              updateArrayLength(1, localMem[1205], 1);
              ip = 2700;
      end

       2700 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 1] = heapMem[localMem[1205]*6 + 1];
              updateArrayLength(1, localMem[1210], 1);
              ip = 2701;
      end

       2701 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1213] = !heapMem[localMem[1202]*6 + 6];
              ip = 2702;
      end

       2702 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1213] != 0 ? 2731 : 2703;
      end

       2703 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1214] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1214] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1214]] = 0;
              ip = 2704;
      end

       2704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 6] = localMem[1214];
              updateArrayLength(1, localMem[1210], 6);
              ip = 2705;
      end

       2705 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1215] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2706;
      end

       2706 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1216] = heapMem[localMem[1210]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2707;
      end

       2707 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1216] + 0 + i] = heapMem[NArea * localMem[1215] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1216], 0 + i);
                end
              end
              ip = 2708;
      end

       2708 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1217] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2709;
      end

       2709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1218] = heapMem[localMem[1210]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2710;
      end

       2710 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1218] + 0 + i] = heapMem[NArea * localMem[1217] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1218], 0 + i);
                end
              end
              ip = 2711;
      end

       2711 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1219] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2712;
      end

       2712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1220] = heapMem[localMem[1210]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2713;
      end

       2713 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1221] = localMem[1207] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2714;
      end

       2714 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1221]) begin
                  heapMem[NArea * localMem[1220] + 0 + i] = heapMem[NArea * localMem[1219] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1220], 0 + i);
                end
              end
              ip = 2715;
      end

       2715 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1222] = heapMem[localMem[1210]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2716;
      end

       2716 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1223] = localMem[1222] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2717;
      end

       2717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1224] = heapMem[localMem[1210]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2718;
      end

       2718 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2719;
      end

       2719 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1225] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2720;
      end

       2720 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2721;
      end

       2721 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1225] >= localMem[1223] ? 2727 : 2722;
      end

       2722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1226] = heapMem[localMem[1224]*6 + localMem[1225]];
              updateArrayLength(2, 0, 0);
              ip = 2723;
      end

       2723 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1226]*6 + 2] = localMem[1210];
              updateArrayLength(1, localMem[1226], 2);
              ip = 2724;
      end

       2724 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2725;
      end

       2725 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1225] = localMem[1225] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2726;
      end

       2726 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2720;
      end

       2727 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2728;
      end

       2728 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1227] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2729;
      end

       2729 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1227]] = localMem[1208];
              ip = 2730;
      end

       2730 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2738;
      end

       2731 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2732;
      end

       2732 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1228] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2733;
      end

       2733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1229] = heapMem[localMem[1210]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2734;
      end

       2734 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1229] + 0 + i] = heapMem[NArea * localMem[1228] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1229], 0 + i);
                end
              end
              ip = 2735;
      end

       2735 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1230] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2736;
      end

       2736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1231] = heapMem[localMem[1210]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2737;
      end

       2737 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1231] + 0 + i] = heapMem[NArea * localMem[1230] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1231], 0 + i);
                end
              end
              ip = 2738;
      end

       2738 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2739;
      end

       2739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1202]*6 + 0] = localMem[1207];
              updateArrayLength(1, localMem[1202], 0);
              ip = 2740;
      end

       2740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1210]*6 + 2] = localMem[1209];
              updateArrayLength(1, localMem[1210], 2);
              ip = 2741;
      end

       2741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1232] = heapMem[localMem[1209]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2742;
      end

       2742 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1233] = heapMem[localMem[1209]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2743;
      end

       2743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1234] = heapMem[localMem[1233]*6 + localMem[1232]];
              updateArrayLength(2, 0, 0);
              ip = 2744;
      end

       2744 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1234] != localMem[1202] ? 2763 : 2745;
      end

       2745 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1235] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2746;
      end

       2746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1236] = heapMem[localMem[1235]*6 + localMem[1207]];
              updateArrayLength(2, 0, 0);
              ip = 2747;
      end

       2747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1237] = heapMem[localMem[1209]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2748;
      end

       2748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1237]*6 + localMem[1232]] = localMem[1236];
              updateArrayLength(1, localMem[1237], localMem[1232]);
              ip = 2749;
      end

       2749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1238] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2750;
      end

       2750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1239] = heapMem[localMem[1238]*6 + localMem[1207]];
              updateArrayLength(2, 0, 0);
              ip = 2751;
      end

       2751 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1240] = heapMem[localMem[1209]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2752;
      end

       2752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1240]*6 + localMem[1232]] = localMem[1239];
              updateArrayLength(1, localMem[1240], localMem[1232]);
              ip = 2753;
      end

       2753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1241] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2754;
      end

       2754 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1241]] = localMem[1207];
              ip = 2755;
      end

       2755 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1242] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2756;
      end

       2756 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1242]] = localMem[1207];
              ip = 2757;
      end

       2757 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1243] = localMem[1232] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2758;
      end

       2758 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1209]*6 + 0] = localMem[1243];
              updateArrayLength(1, localMem[1209], 0);
              ip = 2759;
      end

       2759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1244] = heapMem[localMem[1209]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2760;
      end

       2760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1244]*6 + localMem[1243]] = localMem[1210];
              updateArrayLength(1, localMem[1244], localMem[1243]);
              ip = 2761;
      end

       2761 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2901;
      end

       2762 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2785;
      end

       2763 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2764;
      end

       2764 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 2765;
      end

       2765 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1245] = heapMem[localMem[1209]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2766;
      end

       2766 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1246] = 0; k = arraySizes[localMem[1245]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1245] * NArea + i] == localMem[1202]) localMem[1246] = i + 1;
              end
              ip = 2767;
      end

       2767 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1246] = localMem[1246] - 1;
              updateArrayLength(2, 0, 0);
              ip = 2768;
      end

       2768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1247] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2769;
      end

       2769 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1248] = heapMem[localMem[1247]*6 + localMem[1207]];
              updateArrayLength(2, 0, 0);
              ip = 2770;
      end

       2770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1249] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2771;
      end

       2771 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1250] = heapMem[localMem[1249]*6 + localMem[1207]];
              updateArrayLength(2, 0, 0);
              ip = 2772;
      end

       2772 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1251] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2773;
      end

       2773 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1251]] = localMem[1207];
              ip = 2774;
      end

       2774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1252] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2775;
      end

       2775 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1252]] = localMem[1207];
              ip = 2776;
      end

       2776 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1253] = heapMem[localMem[1209]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2777;
      end

       2777 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1253] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1246], localMem[1253], arraySizes[localMem[1253]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1246] && i <= arraySizes[localMem[1253]]) begin
                  heapMem[NArea * localMem[1253] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1253] + localMem[1246]] = localMem[1248];                                    // Insert new value
              arraySizes[localMem[1253]] = arraySizes[localMem[1253]] + 1;                              // Increase array size
              ip = 2778;
      end

       2778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1254] = heapMem[localMem[1209]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2779;
      end

       2779 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1254] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1246], localMem[1254], arraySizes[localMem[1254]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1246] && i <= arraySizes[localMem[1254]]) begin
                  heapMem[NArea * localMem[1254] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1254] + localMem[1246]] = localMem[1250];                                    // Insert new value
              arraySizes[localMem[1254]] = arraySizes[localMem[1254]] + 1;                              // Increase array size
              ip = 2780;
      end

       2780 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1255] = heapMem[localMem[1209]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2781;
      end

       2781 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1256] = localMem[1246] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2782;
      end

       2782 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1255] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1256], localMem[1255], arraySizes[localMem[1255]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1256] && i <= arraySizes[localMem[1255]]) begin
                  heapMem[NArea * localMem[1255] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1255] + localMem[1256]] = localMem[1210];                                    // Insert new value
              arraySizes[localMem[1255]] = arraySizes[localMem[1255]] + 1;                              // Increase array size
              ip = 2783;
      end

       2783 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1209]*6 + 0] = heapMem[localMem[1209]*6 + 0] + 1;
              updateArrayLength(1, localMem[1209], 0);
              ip = 2784;
      end

       2784 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2901;
      end

       2785 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2786;
      end

       2786 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2787;
      end

       2787 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1257] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1257] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1257]] = 0;
              ip = 2788;
      end

       2788 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 0] = localMem[1207];
              updateArrayLength(1, localMem[1257], 0);
              ip = 2789;
      end

       2789 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 2] = 0;
              updateArrayLength(1, localMem[1257], 2);
              ip = 2790;
      end

       2790 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1258] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1258] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1258]] = 0;
              ip = 2791;
      end

       2791 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 4] = localMem[1258];
              updateArrayLength(1, localMem[1257], 4);
              ip = 2792;
      end

       2792 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1259] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1259] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1259]] = 0;
              ip = 2793;
      end

       2793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 5] = localMem[1259];
              updateArrayLength(1, localMem[1257], 5);
              ip = 2794;
      end

       2794 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 6] = 0;
              updateArrayLength(1, localMem[1257], 6);
              ip = 2795;
      end

       2795 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 3] = localMem[1205];
              updateArrayLength(1, localMem[1257], 3);
              ip = 2796;
      end

       2796 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1205]*6 + 1] = heapMem[localMem[1205]*6 + 1] + 1;
              updateArrayLength(1, localMem[1205], 1);
              ip = 2797;
      end

       2797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 1] = heapMem[localMem[1205]*6 + 1];
              updateArrayLength(1, localMem[1257], 1);
              ip = 2798;
      end

       2798 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1260] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1260] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1260]] = 0;
              ip = 2799;
      end

       2799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 0] = localMem[1207];
              updateArrayLength(1, localMem[1260], 0);
              ip = 2800;
      end

       2800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 2] = 0;
              updateArrayLength(1, localMem[1260], 2);
              ip = 2801;
      end

       2801 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1261] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1261] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1261]] = 0;
              ip = 2802;
      end

       2802 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 4] = localMem[1261];
              updateArrayLength(1, localMem[1260], 4);
              ip = 2803;
      end

       2803 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1262] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1262] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1262]] = 0;
              ip = 2804;
      end

       2804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 5] = localMem[1262];
              updateArrayLength(1, localMem[1260], 5);
              ip = 2805;
      end

       2805 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 6] = 0;
              updateArrayLength(1, localMem[1260], 6);
              ip = 2806;
      end

       2806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 3] = localMem[1205];
              updateArrayLength(1, localMem[1260], 3);
              ip = 2807;
      end

       2807 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1205]*6 + 1] = heapMem[localMem[1205]*6 + 1] + 1;
              updateArrayLength(1, localMem[1205], 1);
              ip = 2808;
      end

       2808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 1] = heapMem[localMem[1205]*6 + 1];
              updateArrayLength(1, localMem[1260], 1);
              ip = 2809;
      end

       2809 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1263] = !heapMem[localMem[1202]*6 + 6];
              ip = 2810;
      end

       2810 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1263] != 0 ? 2862 : 2811;
      end

       2811 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1264] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1264] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1264]] = 0;
              ip = 2812;
      end

       2812 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 6] = localMem[1264];
              updateArrayLength(1, localMem[1257], 6);
              ip = 2813;
      end

       2813 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1265] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1265] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1265]] = 0;
              ip = 2814;
      end

       2814 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 6] = localMem[1265];
              updateArrayLength(1, localMem[1260], 6);
              ip = 2815;
      end

       2815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1266] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2816;
      end

       2816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1267] = heapMem[localMem[1257]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2817;
      end

       2817 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1267] + 0 + i] = heapMem[NArea * localMem[1266] + 0 + i];
                  updateArrayLength(1, localMem[1267], 0 + i);
                end
              end
              ip = 2818;
      end

       2818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1268] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2819;
      end

       2819 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1269] = heapMem[localMem[1257]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2820;
      end

       2820 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1269] + 0 + i] = heapMem[NArea * localMem[1268] + 0 + i];
                  updateArrayLength(1, localMem[1269], 0 + i);
                end
              end
              ip = 2821;
      end

       2821 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1270] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2822;
      end

       2822 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1271] = heapMem[localMem[1257]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2823;
      end

       2823 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1272] = localMem[1207] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2824;
      end

       2824 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1272]) begin
                  heapMem[NArea * localMem[1271] + 0 + i] = heapMem[NArea * localMem[1270] + 0 + i];
                  updateArrayLength(1, localMem[1271], 0 + i);
                end
              end
              ip = 2825;
      end

       2825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1273] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2826;
      end

       2826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1274] = heapMem[localMem[1260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2827;
      end

       2827 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1274] + 0 + i] = heapMem[NArea * localMem[1273] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1274], 0 + i);
                end
              end
              ip = 2828;
      end

       2828 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1275] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2829;
      end

       2829 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1276] = heapMem[localMem[1260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2830;
      end

       2830 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1276] + 0 + i] = heapMem[NArea * localMem[1275] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1276], 0 + i);
                end
              end
              ip = 2831;
      end

       2831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1277] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2832;
      end

       2832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1278] = heapMem[localMem[1260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2833;
      end

       2833 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1279] = localMem[1207] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2834;
      end

       2834 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1279]) begin
                  heapMem[NArea * localMem[1278] + 0 + i] = heapMem[NArea * localMem[1277] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1278], 0 + i);
                end
              end
              ip = 2835;
      end

       2835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1280] = heapMem[localMem[1257]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2836;
      end

       2836 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1281] = localMem[1280] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2837;
      end

       2837 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1282] = heapMem[localMem[1257]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2838;
      end

       2838 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2839;
      end

       2839 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1283] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2840;
      end

       2840 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2841;
      end

       2841 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1283] >= localMem[1281] ? 2847 : 2842;
      end

       2842 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1284] = heapMem[localMem[1282]*6 + localMem[1283]];
              updateArrayLength(2, 0, 0);
              ip = 2843;
      end

       2843 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1284]*6 + 2] = localMem[1257];
              updateArrayLength(1, localMem[1284], 2);
              ip = 2844;
      end

       2844 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2845;
      end

       2845 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1283] = localMem[1283] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2846;
      end

       2846 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2840;
      end

       2847 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2848;
      end

       2848 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1285] = heapMem[localMem[1260]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2849;
      end

       2849 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1286] = localMem[1285] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2850;
      end

       2850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1287] = heapMem[localMem[1260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2851;
      end

       2851 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2852;
      end

       2852 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1288] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2853;
      end

       2853 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2854;
      end

       2854 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1288] >= localMem[1286] ? 2860 : 2855;
      end

       2855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1289] = heapMem[localMem[1287]*6 + localMem[1288]];
              updateArrayLength(2, 0, 0);
              ip = 2856;
      end

       2856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1289]*6 + 2] = localMem[1260];
              updateArrayLength(1, localMem[1289], 2);
              ip = 2857;
      end

       2857 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2858;
      end

       2858 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1288] = localMem[1288] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2859;
      end

       2859 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2853;
      end

       2860 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2861;
      end

       2861 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2877;
      end

       2862 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2863;
      end

       2863 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1290] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1290] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1290]] = 0;
              ip = 2864;
      end

       2864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1202]*6 + 6] = localMem[1290];
              updateArrayLength(1, localMem[1202], 6);
              ip = 2865;
      end

       2865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1291] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2866;
      end

       2866 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1292] = heapMem[localMem[1257]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2867;
      end

       2867 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1292] + 0 + i] = heapMem[NArea * localMem[1291] + 0 + i];
                  updateArrayLength(1, localMem[1292], 0 + i);
                end
              end
              ip = 2868;
      end

       2868 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1293] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2869;
      end

       2869 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1294] = heapMem[localMem[1257]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2870;
      end

       2870 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1294] + 0 + i] = heapMem[NArea * localMem[1293] + 0 + i];
                  updateArrayLength(1, localMem[1294], 0 + i);
                end
              end
              ip = 2871;
      end

       2871 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1295] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2872;
      end

       2872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1296] = heapMem[localMem[1260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2873;
      end

       2873 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1296] + 0 + i] = heapMem[NArea * localMem[1295] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1296], 0 + i);
                end
              end
              ip = 2874;
      end

       2874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1297] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2875;
      end

       2875 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1298] = heapMem[localMem[1260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2876;
      end

       2876 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1207]) begin
                  heapMem[NArea * localMem[1298] + 0 + i] = heapMem[NArea * localMem[1297] + localMem[1208] + i];
                  updateArrayLength(1, localMem[1298], 0 + i);
                end
              end
              ip = 2877;
      end

       2877 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2878;
      end

       2878 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1257]*6 + 2] = localMem[1202];
              updateArrayLength(1, localMem[1257], 2);
              ip = 2879;
      end

       2879 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1260]*6 + 2] = localMem[1202];
              updateArrayLength(1, localMem[1260], 2);
              ip = 2880;
      end

       2880 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1299] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2881;
      end

       2881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1300] = heapMem[localMem[1299]*6 + localMem[1207]];
              updateArrayLength(2, 0, 0);
              ip = 2882;
      end

       2882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1301] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2883;
      end

       2883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1302] = heapMem[localMem[1301]*6 + localMem[1207]];
              updateArrayLength(2, 0, 0);
              ip = 2884;
      end

       2884 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1303] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2885;
      end

       2885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1303]*6 + 0] = localMem[1300];
              updateArrayLength(1, localMem[1303], 0);
              ip = 2886;
      end

       2886 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1304] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2887;
      end

       2887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1304]*6 + 0] = localMem[1302];
              updateArrayLength(1, localMem[1304], 0);
              ip = 2888;
      end

       2888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1305] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2889;
      end

       2889 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1305]*6 + 0] = localMem[1257];
              updateArrayLength(1, localMem[1305], 0);
              ip = 2890;
      end

       2890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1306] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2891;
      end

       2891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1306]*6 + 1] = localMem[1260];
              updateArrayLength(1, localMem[1306], 1);
              ip = 2892;
      end

       2892 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1202]*6 + 0] = 1;
              updateArrayLength(1, localMem[1202], 0);
              ip = 2893;
      end

       2893 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1307] = heapMem[localMem[1202]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2894;
      end

       2894 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1307]] = 1;
              ip = 2895;
      end

       2895 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1308] = heapMem[localMem[1202]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2896;
      end

       2896 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1308]] = 1;
              ip = 2897;
      end

       2897 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1309] = heapMem[localMem[1202]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2898;
      end

       2898 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1309]] = 2;
              ip = 2899;
      end

       2899 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2901;
      end

       2900 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2906;
      end

       2901 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2902;
      end

       2902 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1203] = 1;
              updateArrayLength(2, 0, 0);
              ip = 2903;
      end

       2903 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2906;
      end

       2904 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2905;
      end

       2905 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1203] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2906;
      end

       2906 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2907;
      end

       2907 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1203] != 0 ? 2909 : 2908;
      end

       2908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[974] = localMem[1202];
              updateArrayLength(2, 0, 0);
              ip = 2909;
      end

       2909 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2910;
      end

       2910 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2911;
      end

       2911 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1082] = localMem[1082] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2912;
      end

       2912 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2414;
      end

       2913 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2914;
      end

       2914 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
            ip = 2915;
      end

       2915 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2916;
      end

       2916 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2917;
      end

       2917 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2918;
      end

       2918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1310] = heapMem[localMem[951]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2919;
      end

       2919 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1311] = heapMem[localMem[951]*6 + 1];
              updateArrayLength(2, 0, 0);
              ip = 2920;
      end

       2920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1312] = heapMem[localMem[951]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2921;
      end

       2921 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1311] != 1 ? 2925 : 2922;
      end

       2922 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1313] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2923;
      end

       2923 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1313]*6 + localMem[1312]] = 33;
              updateArrayLength(1, localMem[1313], localMem[1312]);
              ip = 2924;
      end

       2924 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3171;
      end

       2925 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2926;
      end

       2926 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1311] != 2 ? 2934 : 2927;
      end

       2927 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1314] = localMem[1312] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2928;
      end

       2928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1315] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2929;
      end

       2929 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1315] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1314], localMem[1315], arraySizes[localMem[1315]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1314] && i <= arraySizes[localMem[1315]]) begin
                  heapMem[NArea * localMem[1315] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1315] + localMem[1314]] = 3;                                    // Insert new value
              arraySizes[localMem[1315]] = arraySizes[localMem[1315]] + 1;                              // Increase array size
              ip = 2930;
      end

       2930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1316] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2931;
      end

       2931 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1316] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1314], localMem[1316], arraySizes[localMem[1316]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1314] && i <= arraySizes[localMem[1316]]) begin
                  heapMem[NArea * localMem[1316] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1316] + localMem[1314]] = 33;                                    // Insert new value
              arraySizes[localMem[1316]] = arraySizes[localMem[1316]] + 1;                              // Increase array size
              ip = 2932;
      end

       2932 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1310]*6 + 0] = heapMem[localMem[1310]*6 + 0] + 1;
              updateArrayLength(1, localMem[1310], 0);
              ip = 2933;
      end

       2933 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2940;
      end

       2934 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2935;
      end

       2935 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1317] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2936;
      end

       2936 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1317] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1312], localMem[1317], arraySizes[localMem[1317]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1312] && i <= arraySizes[localMem[1317]]) begin
                  heapMem[NArea * localMem[1317] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1317] + localMem[1312]] = 3;                                    // Insert new value
              arraySizes[localMem[1317]] = arraySizes[localMem[1317]] + 1;                              // Increase array size
              ip = 2937;
      end

       2937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1318] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2938;
      end

       2938 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1318] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1312], localMem[1318], arraySizes[localMem[1318]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1312] && i <= arraySizes[localMem[1318]]) begin
                  heapMem[NArea * localMem[1318] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1318] + localMem[1312]] = 33;                                    // Insert new value
              arraySizes[localMem[1318]] = arraySizes[localMem[1318]] + 1;                              // Increase array size
              ip = 2939;
      end

       2939 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1310]*6 + 0] = heapMem[localMem[1310]*6 + 0] + 1;
              updateArrayLength(1, localMem[1310], 0);
              ip = 2940;
      end

       2940 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2941;
      end

       2941 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 2942;
      end

       2942 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2943;
      end

       2943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1320] = heapMem[localMem[1310]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2944;
      end

       2944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1321] = heapMem[localMem[1310]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2945;
      end

       2945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1322] = heapMem[localMem[1321]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2946;
      end

       2946 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1320] <  localMem[1322] ? 3166 : 2947;
      end

       2947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1323] = localMem[1322];
              updateArrayLength(2, 0, 0);
              ip = 2948;
      end

       2948 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1323] = localMem[1323] >> 1;
              ip = 2949;
      end

       2949 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1324] = localMem[1323] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2950;
      end

       2950 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1325] = heapMem[localMem[1310]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2951;
      end

       2951 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1325] == 0 ? 3048 : 2952;
      end

       2952 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1326] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1326] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1326]] = 0;
              ip = 2953;
      end

       2953 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 0] = localMem[1323];
              updateArrayLength(1, localMem[1326], 0);
              ip = 2954;
      end

       2954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 2] = 0;
              updateArrayLength(1, localMem[1326], 2);
              ip = 2955;
      end

       2955 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1327] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1327] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1327]] = 0;
              ip = 2956;
      end

       2956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 4] = localMem[1327];
              updateArrayLength(1, localMem[1326], 4);
              ip = 2957;
      end

       2957 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1328] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1328] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1328]] = 0;
              ip = 2958;
      end

       2958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 5] = localMem[1328];
              updateArrayLength(1, localMem[1326], 5);
              ip = 2959;
      end

       2959 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 6] = 0;
              updateArrayLength(1, localMem[1326], 6);
              ip = 2960;
      end

       2960 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 3] = localMem[1321];
              updateArrayLength(1, localMem[1326], 3);
              ip = 2961;
      end

       2961 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1321]*6 + 1] = heapMem[localMem[1321]*6 + 1] + 1;
              updateArrayLength(1, localMem[1321], 1);
              ip = 2962;
      end

       2962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 1] = heapMem[localMem[1321]*6 + 1];
              updateArrayLength(1, localMem[1326], 1);
              ip = 2963;
      end

       2963 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1329] = !heapMem[localMem[1310]*6 + 6];
              ip = 2964;
      end

       2964 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1329] != 0 ? 2993 : 2965;
      end

       2965 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1330] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1330] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1330]] = 0;
              ip = 2966;
      end

       2966 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 6] = localMem[1330];
              updateArrayLength(1, localMem[1326], 6);
              ip = 2967;
      end

       2967 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1331] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2968;
      end

       2968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1332] = heapMem[localMem[1326]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2969;
      end

       2969 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1332] + 0 + i] = heapMem[NArea * localMem[1331] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1332], 0 + i);
                end
              end
              ip = 2970;
      end

       2970 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1333] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2971;
      end

       2971 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1334] = heapMem[localMem[1326]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2972;
      end

       2972 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1334] + 0 + i] = heapMem[NArea * localMem[1333] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1334], 0 + i);
                end
              end
              ip = 2973;
      end

       2973 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1335] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2974;
      end

       2974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1336] = heapMem[localMem[1326]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2975;
      end

       2975 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1337] = localMem[1323] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2976;
      end

       2976 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1337]) begin
                  heapMem[NArea * localMem[1336] + 0 + i] = heapMem[NArea * localMem[1335] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1336], 0 + i);
                end
              end
              ip = 2977;
      end

       2977 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1338] = heapMem[localMem[1326]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2978;
      end

       2978 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1339] = localMem[1338] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2979;
      end

       2979 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1340] = heapMem[localMem[1326]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2980;
      end

       2980 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2981;
      end

       2981 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1341] = 0;
              updateArrayLength(2, 0, 0);
              ip = 2982;
      end

       2982 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2983;
      end

       2983 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1341] >= localMem[1339] ? 2989 : 2984;
      end

       2984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1342] = heapMem[localMem[1340]*6 + localMem[1341]];
              updateArrayLength(2, 0, 0);
              ip = 2985;
      end

       2985 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1342]*6 + 2] = localMem[1326];
              updateArrayLength(1, localMem[1342], 2);
              ip = 2986;
      end

       2986 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2987;
      end

       2987 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1341] = localMem[1341] + 1;
              updateArrayLength(2, 0, 0);
              ip = 2988;
      end

       2988 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2982;
      end

       2989 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2990;
      end

       2990 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1343] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 2991;
      end

       2991 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1343]] = localMem[1324];
              ip = 2992;
      end

       2992 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3000;
      end

       2993 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2994;
      end

       2994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1344] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2995;
      end

       2995 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1345] = heapMem[localMem[1326]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2996;
      end

       2996 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1345] + 0 + i] = heapMem[NArea * localMem[1344] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1345], 0 + i);
                end
              end
              ip = 2997;
      end

       2997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1346] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2998;
      end

       2998 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1347] = heapMem[localMem[1326]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2999;
      end

       2999 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1347] + 0 + i] = heapMem[NArea * localMem[1346] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1347], 0 + i);
                end
              end
              ip = 3000;
      end

       3000 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3001;
      end

       3001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1310]*6 + 0] = localMem[1323];
              updateArrayLength(1, localMem[1310], 0);
              ip = 3002;
      end

       3002 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1326]*6 + 2] = localMem[1325];
              updateArrayLength(1, localMem[1326], 2);
              ip = 3003;
      end

       3003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1348] = heapMem[localMem[1325]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3004;
      end

       3004 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1349] = heapMem[localMem[1325]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3005;
      end

       3005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1350] = heapMem[localMem[1349]*6 + localMem[1348]];
              updateArrayLength(2, 0, 0);
              ip = 3006;
      end

       3006 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1350] != localMem[1310] ? 3025 : 3007;
      end

       3007 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1351] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3008;
      end

       3008 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1352] = heapMem[localMem[1351]*6 + localMem[1323]];
              updateArrayLength(2, 0, 0);
              ip = 3009;
      end

       3009 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1353] = heapMem[localMem[1325]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3010;
      end

       3010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1353]*6 + localMem[1348]] = localMem[1352];
              updateArrayLength(1, localMem[1353], localMem[1348]);
              ip = 3011;
      end

       3011 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1354] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3012;
      end

       3012 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1355] = heapMem[localMem[1354]*6 + localMem[1323]];
              updateArrayLength(2, 0, 0);
              ip = 3013;
      end

       3013 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1356] = heapMem[localMem[1325]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3014;
      end

       3014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1356]*6 + localMem[1348]] = localMem[1355];
              updateArrayLength(1, localMem[1356], localMem[1348]);
              ip = 3015;
      end

       3015 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1357] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3016;
      end

       3016 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1357]] = localMem[1323];
              ip = 3017;
      end

       3017 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1358] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3018;
      end

       3018 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1358]] = localMem[1323];
              ip = 3019;
      end

       3019 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1359] = localMem[1348] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3020;
      end

       3020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1325]*6 + 0] = localMem[1359];
              updateArrayLength(1, localMem[1325], 0);
              ip = 3021;
      end

       3021 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1360] = heapMem[localMem[1325]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3022;
      end

       3022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1360]*6 + localMem[1359]] = localMem[1326];
              updateArrayLength(1, localMem[1360], localMem[1359]);
              ip = 3023;
      end

       3023 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3163;
      end

       3024 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3047;
      end

       3025 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3026;
      end

       3026 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 3027;
      end

       3027 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1361] = heapMem[localMem[1325]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3028;
      end

       3028 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1362] = 0; k = arraySizes[localMem[1361]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1361] * NArea + i] == localMem[1310]) localMem[1362] = i + 1;
              end
              ip = 3029;
      end

       3029 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1362] = localMem[1362] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3030;
      end

       3030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1363] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3031;
      end

       3031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1364] = heapMem[localMem[1363]*6 + localMem[1323]];
              updateArrayLength(2, 0, 0);
              ip = 3032;
      end

       3032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1365] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3033;
      end

       3033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1366] = heapMem[localMem[1365]*6 + localMem[1323]];
              updateArrayLength(2, 0, 0);
              ip = 3034;
      end

       3034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1367] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3035;
      end

       3035 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1367]] = localMem[1323];
              ip = 3036;
      end

       3036 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1368] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3037;
      end

       3037 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1368]] = localMem[1323];
              ip = 3038;
      end

       3038 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1369] = heapMem[localMem[1325]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3039;
      end

       3039 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1369] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1362], localMem[1369], arraySizes[localMem[1369]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1362] && i <= arraySizes[localMem[1369]]) begin
                  heapMem[NArea * localMem[1369] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1369] + localMem[1362]] = localMem[1364];                                    // Insert new value
              arraySizes[localMem[1369]] = arraySizes[localMem[1369]] + 1;                              // Increase array size
              ip = 3040;
      end

       3040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1370] = heapMem[localMem[1325]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3041;
      end

       3041 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1370] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1362], localMem[1370], arraySizes[localMem[1370]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1362] && i <= arraySizes[localMem[1370]]) begin
                  heapMem[NArea * localMem[1370] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1370] + localMem[1362]] = localMem[1366];                                    // Insert new value
              arraySizes[localMem[1370]] = arraySizes[localMem[1370]] + 1;                              // Increase array size
              ip = 3042;
      end

       3042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1371] = heapMem[localMem[1325]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3043;
      end

       3043 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1372] = localMem[1362] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3044;
      end

       3044 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1371] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1372], localMem[1371], arraySizes[localMem[1371]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1372] && i <= arraySizes[localMem[1371]]) begin
                  heapMem[NArea * localMem[1371] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1371] + localMem[1372]] = localMem[1326];                                    // Insert new value
              arraySizes[localMem[1371]] = arraySizes[localMem[1371]] + 1;                              // Increase array size
              ip = 3045;
      end

       3045 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1325]*6 + 0] = heapMem[localMem[1325]*6 + 0] + 1;
              updateArrayLength(1, localMem[1325], 0);
              ip = 3046;
      end

       3046 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3163;
      end

       3047 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3048;
      end

       3048 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3049;
      end

       3049 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1373] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1373] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1373]] = 0;
              ip = 3050;
      end

       3050 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 0] = localMem[1323];
              updateArrayLength(1, localMem[1373], 0);
              ip = 3051;
      end

       3051 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 2] = 0;
              updateArrayLength(1, localMem[1373], 2);
              ip = 3052;
      end

       3052 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1374] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1374] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1374]] = 0;
              ip = 3053;
      end

       3053 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 4] = localMem[1374];
              updateArrayLength(1, localMem[1373], 4);
              ip = 3054;
      end

       3054 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1375] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1375] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1375]] = 0;
              ip = 3055;
      end

       3055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 5] = localMem[1375];
              updateArrayLength(1, localMem[1373], 5);
              ip = 3056;
      end

       3056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 6] = 0;
              updateArrayLength(1, localMem[1373], 6);
              ip = 3057;
      end

       3057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 3] = localMem[1321];
              updateArrayLength(1, localMem[1373], 3);
              ip = 3058;
      end

       3058 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1321]*6 + 1] = heapMem[localMem[1321]*6 + 1] + 1;
              updateArrayLength(1, localMem[1321], 1);
              ip = 3059;
      end

       3059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 1] = heapMem[localMem[1321]*6 + 1];
              updateArrayLength(1, localMem[1373], 1);
              ip = 3060;
      end

       3060 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1376] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1376] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1376]] = 0;
              ip = 3061;
      end

       3061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 0] = localMem[1323];
              updateArrayLength(1, localMem[1376], 0);
              ip = 3062;
      end

       3062 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 2] = 0;
              updateArrayLength(1, localMem[1376], 2);
              ip = 3063;
      end

       3063 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1377] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1377] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1377]] = 0;
              ip = 3064;
      end

       3064 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 4] = localMem[1377];
              updateArrayLength(1, localMem[1376], 4);
              ip = 3065;
      end

       3065 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1378] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1378] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1378]] = 0;
              ip = 3066;
      end

       3066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 5] = localMem[1378];
              updateArrayLength(1, localMem[1376], 5);
              ip = 3067;
      end

       3067 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 6] = 0;
              updateArrayLength(1, localMem[1376], 6);
              ip = 3068;
      end

       3068 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 3] = localMem[1321];
              updateArrayLength(1, localMem[1376], 3);
              ip = 3069;
      end

       3069 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1321]*6 + 1] = heapMem[localMem[1321]*6 + 1] + 1;
              updateArrayLength(1, localMem[1321], 1);
              ip = 3070;
      end

       3070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 1] = heapMem[localMem[1321]*6 + 1];
              updateArrayLength(1, localMem[1376], 1);
              ip = 3071;
      end

       3071 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1379] = !heapMem[localMem[1310]*6 + 6];
              ip = 3072;
      end

       3072 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1379] != 0 ? 3124 : 3073;
      end

       3073 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1380] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1380] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1380]] = 0;
              ip = 3074;
      end

       3074 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 6] = localMem[1380];
              updateArrayLength(1, localMem[1373], 6);
              ip = 3075;
      end

       3075 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1381] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1381] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1381]] = 0;
              ip = 3076;
      end

       3076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 6] = localMem[1381];
              updateArrayLength(1, localMem[1376], 6);
              ip = 3077;
      end

       3077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1382] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3078;
      end

       3078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1383] = heapMem[localMem[1373]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3079;
      end

       3079 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1383] + 0 + i] = heapMem[NArea * localMem[1382] + 0 + i];
                  updateArrayLength(1, localMem[1383], 0 + i);
                end
              end
              ip = 3080;
      end

       3080 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1384] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3081;
      end

       3081 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1385] = heapMem[localMem[1373]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3082;
      end

       3082 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1385] + 0 + i] = heapMem[NArea * localMem[1384] + 0 + i];
                  updateArrayLength(1, localMem[1385], 0 + i);
                end
              end
              ip = 3083;
      end

       3083 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1386] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3084;
      end

       3084 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1387] = heapMem[localMem[1373]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3085;
      end

       3085 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1388] = localMem[1323] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3086;
      end

       3086 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1388]) begin
                  heapMem[NArea * localMem[1387] + 0 + i] = heapMem[NArea * localMem[1386] + 0 + i];
                  updateArrayLength(1, localMem[1387], 0 + i);
                end
              end
              ip = 3087;
      end

       3087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1389] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3088;
      end

       3088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1390] = heapMem[localMem[1376]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3089;
      end

       3089 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1390] + 0 + i] = heapMem[NArea * localMem[1389] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1390], 0 + i);
                end
              end
              ip = 3090;
      end

       3090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1391] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3091;
      end

       3091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1392] = heapMem[localMem[1376]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3092;
      end

       3092 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1392] + 0 + i] = heapMem[NArea * localMem[1391] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1392], 0 + i);
                end
              end
              ip = 3093;
      end

       3093 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1393] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3094;
      end

       3094 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1394] = heapMem[localMem[1376]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3095;
      end

       3095 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1395] = localMem[1323] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3096;
      end

       3096 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1395]) begin
                  heapMem[NArea * localMem[1394] + 0 + i] = heapMem[NArea * localMem[1393] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1394], 0 + i);
                end
              end
              ip = 3097;
      end

       3097 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1396] = heapMem[localMem[1373]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3098;
      end

       3098 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1397] = localMem[1396] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3099;
      end

       3099 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1398] = heapMem[localMem[1373]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3100;
      end

       3100 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3101;
      end

       3101 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1399] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3102;
      end

       3102 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3103;
      end

       3103 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1399] >= localMem[1397] ? 3109 : 3104;
      end

       3104 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1400] = heapMem[localMem[1398]*6 + localMem[1399]];
              updateArrayLength(2, 0, 0);
              ip = 3105;
      end

       3105 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1400]*6 + 2] = localMem[1373];
              updateArrayLength(1, localMem[1400], 2);
              ip = 3106;
      end

       3106 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3107;
      end

       3107 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1399] = localMem[1399] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3108;
      end

       3108 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3102;
      end

       3109 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3110;
      end

       3110 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1401] = heapMem[localMem[1376]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3111;
      end

       3111 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1402] = localMem[1401] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3112;
      end

       3112 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1403] = heapMem[localMem[1376]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3113;
      end

       3113 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3114;
      end

       3114 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1404] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3115;
      end

       3115 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3116;
      end

       3116 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1404] >= localMem[1402] ? 3122 : 3117;
      end

       3117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1405] = heapMem[localMem[1403]*6 + localMem[1404]];
              updateArrayLength(2, 0, 0);
              ip = 3118;
      end

       3118 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1405]*6 + 2] = localMem[1376];
              updateArrayLength(1, localMem[1405], 2);
              ip = 3119;
      end

       3119 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3120;
      end

       3120 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1404] = localMem[1404] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3121;
      end

       3121 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3115;
      end

       3122 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3123;
      end

       3123 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3139;
      end

       3124 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3125;
      end

       3125 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1406] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1406] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1406]] = 0;
              ip = 3126;
      end

       3126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1310]*6 + 6] = localMem[1406];
              updateArrayLength(1, localMem[1310], 6);
              ip = 3127;
      end

       3127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1407] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3128;
      end

       3128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1408] = heapMem[localMem[1373]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3129;
      end

       3129 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1408] + 0 + i] = heapMem[NArea * localMem[1407] + 0 + i];
                  updateArrayLength(1, localMem[1408], 0 + i);
                end
              end
              ip = 3130;
      end

       3130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1409] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3131;
      end

       3131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1410] = heapMem[localMem[1373]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3132;
      end

       3132 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1410] + 0 + i] = heapMem[NArea * localMem[1409] + 0 + i];
                  updateArrayLength(1, localMem[1410], 0 + i);
                end
              end
              ip = 3133;
      end

       3133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1411] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3134;
      end

       3134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1412] = heapMem[localMem[1376]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3135;
      end

       3135 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1412] + 0 + i] = heapMem[NArea * localMem[1411] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1412], 0 + i);
                end
              end
              ip = 3136;
      end

       3136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1413] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3137;
      end

       3137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1414] = heapMem[localMem[1376]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3138;
      end

       3138 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1323]) begin
                  heapMem[NArea * localMem[1414] + 0 + i] = heapMem[NArea * localMem[1413] + localMem[1324] + i];
                  updateArrayLength(1, localMem[1414], 0 + i);
                end
              end
              ip = 3139;
      end

       3139 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3140;
      end

       3140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1373]*6 + 2] = localMem[1310];
              updateArrayLength(1, localMem[1373], 2);
              ip = 3141;
      end

       3141 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1376]*6 + 2] = localMem[1310];
              updateArrayLength(1, localMem[1376], 2);
              ip = 3142;
      end

       3142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1415] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3143;
      end

       3143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1416] = heapMem[localMem[1415]*6 + localMem[1323]];
              updateArrayLength(2, 0, 0);
              ip = 3144;
      end

       3144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1417] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3145;
      end

       3145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1418] = heapMem[localMem[1417]*6 + localMem[1323]];
              updateArrayLength(2, 0, 0);
              ip = 3146;
      end

       3146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1419] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3147;
      end

       3147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1419]*6 + 0] = localMem[1416];
              updateArrayLength(1, localMem[1419], 0);
              ip = 3148;
      end

       3148 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1420] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3149;
      end

       3149 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1420]*6 + 0] = localMem[1418];
              updateArrayLength(1, localMem[1420], 0);
              ip = 3150;
      end

       3150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1421] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3151;
      end

       3151 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1421]*6 + 0] = localMem[1373];
              updateArrayLength(1, localMem[1421], 0);
              ip = 3152;
      end

       3152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1422] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3153;
      end

       3153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1422]*6 + 1] = localMem[1376];
              updateArrayLength(1, localMem[1422], 1);
              ip = 3154;
      end

       3154 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1310]*6 + 0] = 1;
              updateArrayLength(1, localMem[1310], 0);
              ip = 3155;
      end

       3155 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1423] = heapMem[localMem[1310]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3156;
      end

       3156 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1423]] = 1;
              ip = 3157;
      end

       3157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1424] = heapMem[localMem[1310]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3158;
      end

       3158 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1424]] = 1;
              ip = 3159;
      end

       3159 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1425] = heapMem[localMem[1310]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3160;
      end

       3160 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1425]] = 2;
              ip = 3161;
      end

       3161 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3163;
      end

       3162 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3168;
      end

       3163 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3164;
      end

       3164 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1319] = 1;
              updateArrayLength(2, 0, 0);
              ip = 3165;
      end

       3165 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3168;
      end

       3166 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3167;
      end

       3167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1319] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3168;
      end

       3168 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3169;
      end

       3169 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3170;
      end

       3170 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3171;
      end

       3171 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3172;
      end

       3172 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[951]] = 0;
              freedArrays[freedArraysTop] = localMem[951];
              freedArraysTop = freedArraysTop + 1;
              ip = 3173;
      end

       3173 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1426] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1426] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1426]] = 0;
              ip = 3174;
      end

       3174 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3175;
      end

       3175 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1427] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3176;
      end

       3176 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1427] != 0 ? 3199 : 3177;
      end

       3177 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1428] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1428] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1428]] = 0;
              ip = 3178;
      end

       3178 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 0] = 1;
              updateArrayLength(1, localMem[1428], 0);
              ip = 3179;
      end

       3179 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 2] = 0;
              updateArrayLength(1, localMem[1428], 2);
              ip = 3180;
      end

       3180 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1429] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1429] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1429]] = 0;
              ip = 3181;
      end

       3181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 4] = localMem[1429];
              updateArrayLength(1, localMem[1428], 4);
              ip = 3182;
      end

       3182 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1430] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1430] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1430]] = 0;
              ip = 3183;
      end

       3183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 5] = localMem[1430];
              updateArrayLength(1, localMem[1428], 5);
              ip = 3184;
      end

       3184 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 6] = 0;
              updateArrayLength(1, localMem[1428], 6);
              ip = 3185;
      end

       3185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 3] = localMem[0];
              updateArrayLength(1, localMem[1428], 3);
              ip = 3186;
      end

       3186 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = heapMem[localMem[0]*6 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 3187;
      end

       3187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1428]*6 + 1] = heapMem[localMem[0]*6 + 1];
              updateArrayLength(1, localMem[1428], 1);
              ip = 3188;
      end

       3188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1431] = heapMem[localMem[1428]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3189;
      end

       3189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1431]*6 + 0] = 4;
              updateArrayLength(1, localMem[1431], 0);
              ip = 3190;
      end

       3190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1432] = heapMem[localMem[1428]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3191;
      end

       3191 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1432]*6 + 0] = 44;
              updateArrayLength(1, localMem[1432], 0);
              ip = 3192;
      end

       3192 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 3193;
      end

       3193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = localMem[1428];
              updateArrayLength(1, localMem[0], 3);
              ip = 3194;
      end

       3194 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1433] = heapMem[localMem[1428]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3195;
      end

       3195 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1433]] = 1;
              ip = 3196;
      end

       3196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1434] = heapMem[localMem[1428]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3197;
      end

       3197 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1434]] = 1;
              ip = 3198;
      end

       3198 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4227;
      end

       3199 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3200;
      end

       3200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1435] = heapMem[localMem[1427]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3201;
      end

       3201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1436] = heapMem[localMem[0]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3202;
      end

       3202 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1435] >= localMem[1436] ? 3238 : 3203;
      end

       3203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1437] = heapMem[localMem[1427]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3204;
      end

       3204 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1437] != 0 ? 3237 : 3205;
      end

       3205 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1438] = !heapMem[localMem[1427]*6 + 6];
              ip = 3206;
      end

       3206 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1438] == 0 ? 3236 : 3207;
      end

       3207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1439] = heapMem[localMem[1427]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3208;
      end

       3208 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1440] = 0; k = arraySizes[localMem[1439]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1439] * NArea + i] == 4) localMem[1440] = i + 1;
              end
              ip = 3209;
      end

       3209 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1440] == 0 ? 3214 : 3210;
      end

       3210 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1440] = localMem[1440] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3211;
      end

       3211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1441] = heapMem[localMem[1427]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3212;
      end

       3212 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1441]*6 + localMem[1440]] = 44;
              updateArrayLength(1, localMem[1441], localMem[1440]);
              ip = 3213;
      end

       3213 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4227;
      end

       3214 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3215;
      end

       3215 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1439]] = localMem[1435];
              ip = 3216;
      end

       3216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1442] = heapMem[localMem[1427]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3217;
      end

       3217 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1442]] = localMem[1435];
              ip = 3218;
      end

       3218 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[1439]];
//$display("AAAAA k=%d  source2=%d", k, 4);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[1439] * NArea + i]);
                if (i < k && heapMem[localMem[1439] * NArea + i] > 4) j = j + 1;
              end
              localMem[1443] = j;
              ip = 3219;
      end

       3219 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1443] != 0 ? 3227 : 3220;
      end

       3220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1444] = heapMem[localMem[1427]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3221;
      end

       3221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1444]*6 + localMem[1435]] = 4;
              updateArrayLength(1, localMem[1444], localMem[1435]);
              ip = 3222;
      end

       3222 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1445] = heapMem[localMem[1427]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3223;
      end

       3223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1445]*6 + localMem[1435]] = 44;
              updateArrayLength(1, localMem[1445], localMem[1435]);
              ip = 3224;
      end

       3224 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1427]*6 + 0] = localMem[1435] + 1;
              updateArrayLength(1, localMem[1427], 0);
              ip = 3225;
      end

       3225 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 3226;
      end

       3226 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4227;
      end

       3227 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3228;
      end

       3228 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[1439]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1439] * NArea + i] < 4) j = j + 1;
              end
              localMem[1446] = j;
              ip = 3229;
      end

       3229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1447] = heapMem[localMem[1427]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3230;
      end

       3230 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1447] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1446], localMem[1447], arraySizes[localMem[1447]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1446] && i <= arraySizes[localMem[1447]]) begin
                  heapMem[NArea * localMem[1447] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1447] + localMem[1446]] = 4;                                    // Insert new value
              arraySizes[localMem[1447]] = arraySizes[localMem[1447]] + 1;                              // Increase array size
              ip = 3231;
      end

       3231 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1448] = heapMem[localMem[1427]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3232;
      end

       3232 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1448] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1446], localMem[1448], arraySizes[localMem[1448]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1446] && i <= arraySizes[localMem[1448]]) begin
                  heapMem[NArea * localMem[1448] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1448] + localMem[1446]] = 44;                                    // Insert new value
              arraySizes[localMem[1448]] = arraySizes[localMem[1448]] + 1;                              // Increase array size
              ip = 3233;
      end

       3233 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1427]*6 + 0] = heapMem[localMem[1427]*6 + 0] + 1;
              updateArrayLength(1, localMem[1427], 0);
              ip = 3234;
      end

       3234 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 3235;
      end

       3235 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4227;
      end

       3236 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3237;
      end

       3237 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3238;
      end

       3238 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3239;
      end

       3239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1449] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3240;
      end

       3240 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3241;
      end

       3241 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1451] = heapMem[localMem[1449]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3242;
      end

       3242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1452] = heapMem[localMem[1449]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3243;
      end

       3243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1453] = heapMem[localMem[1452]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3244;
      end

       3244 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1451] <  localMem[1453] ? 3464 : 3245;
      end

       3245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1454] = localMem[1453];
              updateArrayLength(2, 0, 0);
              ip = 3246;
      end

       3246 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1454] = localMem[1454] >> 1;
              ip = 3247;
      end

       3247 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1455] = localMem[1454] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3248;
      end

       3248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1456] = heapMem[localMem[1449]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3249;
      end

       3249 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1456] == 0 ? 3346 : 3250;
      end

       3250 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1457] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1457] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1457]] = 0;
              ip = 3251;
      end

       3251 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 0] = localMem[1454];
              updateArrayLength(1, localMem[1457], 0);
              ip = 3252;
      end

       3252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 2] = 0;
              updateArrayLength(1, localMem[1457], 2);
              ip = 3253;
      end

       3253 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1458] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1458] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1458]] = 0;
              ip = 3254;
      end

       3254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 4] = localMem[1458];
              updateArrayLength(1, localMem[1457], 4);
              ip = 3255;
      end

       3255 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1459] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1459] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1459]] = 0;
              ip = 3256;
      end

       3256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 5] = localMem[1459];
              updateArrayLength(1, localMem[1457], 5);
              ip = 3257;
      end

       3257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 6] = 0;
              updateArrayLength(1, localMem[1457], 6);
              ip = 3258;
      end

       3258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 3] = localMem[1452];
              updateArrayLength(1, localMem[1457], 3);
              ip = 3259;
      end

       3259 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1452]*6 + 1] = heapMem[localMem[1452]*6 + 1] + 1;
              updateArrayLength(1, localMem[1452], 1);
              ip = 3260;
      end

       3260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 1] = heapMem[localMem[1452]*6 + 1];
              updateArrayLength(1, localMem[1457], 1);
              ip = 3261;
      end

       3261 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1460] = !heapMem[localMem[1449]*6 + 6];
              ip = 3262;
      end

       3262 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1460] != 0 ? 3291 : 3263;
      end

       3263 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1461] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1461] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1461]] = 0;
              ip = 3264;
      end

       3264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 6] = localMem[1461];
              updateArrayLength(1, localMem[1457], 6);
              ip = 3265;
      end

       3265 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1462] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3266;
      end

       3266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1463] = heapMem[localMem[1457]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3267;
      end

       3267 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1463] + 0 + i] = heapMem[NArea * localMem[1462] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1463], 0 + i);
                end
              end
              ip = 3268;
      end

       3268 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1464] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3269;
      end

       3269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1465] = heapMem[localMem[1457]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3270;
      end

       3270 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1465] + 0 + i] = heapMem[NArea * localMem[1464] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1465], 0 + i);
                end
              end
              ip = 3271;
      end

       3271 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1466] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3272;
      end

       3272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1467] = heapMem[localMem[1457]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3273;
      end

       3273 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1468] = localMem[1454] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3274;
      end

       3274 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1468]) begin
                  heapMem[NArea * localMem[1467] + 0 + i] = heapMem[NArea * localMem[1466] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1467], 0 + i);
                end
              end
              ip = 3275;
      end

       3275 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1469] = heapMem[localMem[1457]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3276;
      end

       3276 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1470] = localMem[1469] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3277;
      end

       3277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1471] = heapMem[localMem[1457]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3278;
      end

       3278 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3279;
      end

       3279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1472] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3280;
      end

       3280 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3281;
      end

       3281 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1472] >= localMem[1470] ? 3287 : 3282;
      end

       3282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1473] = heapMem[localMem[1471]*6 + localMem[1472]];
              updateArrayLength(2, 0, 0);
              ip = 3283;
      end

       3283 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1473]*6 + 2] = localMem[1457];
              updateArrayLength(1, localMem[1473], 2);
              ip = 3284;
      end

       3284 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3285;
      end

       3285 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1472] = localMem[1472] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3286;
      end

       3286 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3280;
      end

       3287 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3288;
      end

       3288 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1474] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3289;
      end

       3289 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1474]] = localMem[1455];
              ip = 3290;
      end

       3290 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3298;
      end

       3291 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3292;
      end

       3292 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1475] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3293;
      end

       3293 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1476] = heapMem[localMem[1457]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3294;
      end

       3294 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1476] + 0 + i] = heapMem[NArea * localMem[1475] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1476], 0 + i);
                end
              end
              ip = 3295;
      end

       3295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1477] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3296;
      end

       3296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1478] = heapMem[localMem[1457]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3297;
      end

       3297 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1478] + 0 + i] = heapMem[NArea * localMem[1477] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1478], 0 + i);
                end
              end
              ip = 3298;
      end

       3298 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3299;
      end

       3299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1449]*6 + 0] = localMem[1454];
              updateArrayLength(1, localMem[1449], 0);
              ip = 3300;
      end

       3300 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1457]*6 + 2] = localMem[1456];
              updateArrayLength(1, localMem[1457], 2);
              ip = 3301;
      end

       3301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1479] = heapMem[localMem[1456]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3302;
      end

       3302 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1480] = heapMem[localMem[1456]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3303;
      end

       3303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1481] = heapMem[localMem[1480]*6 + localMem[1479]];
              updateArrayLength(2, 0, 0);
              ip = 3304;
      end

       3304 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1481] != localMem[1449] ? 3323 : 3305;
      end

       3305 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1482] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3306;
      end

       3306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1483] = heapMem[localMem[1482]*6 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3307;
      end

       3307 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1484] = heapMem[localMem[1456]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3308;
      end

       3308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1484]*6 + localMem[1479]] = localMem[1483];
              updateArrayLength(1, localMem[1484], localMem[1479]);
              ip = 3309;
      end

       3309 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1485] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3310;
      end

       3310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1486] = heapMem[localMem[1485]*6 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3311;
      end

       3311 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1487] = heapMem[localMem[1456]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3312;
      end

       3312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1487]*6 + localMem[1479]] = localMem[1486];
              updateArrayLength(1, localMem[1487], localMem[1479]);
              ip = 3313;
      end

       3313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1488] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3314;
      end

       3314 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1488]] = localMem[1454];
              ip = 3315;
      end

       3315 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1489] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3316;
      end

       3316 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1489]] = localMem[1454];
              ip = 3317;
      end

       3317 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1490] = localMem[1479] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3318;
      end

       3318 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1456]*6 + 0] = localMem[1490];
              updateArrayLength(1, localMem[1456], 0);
              ip = 3319;
      end

       3319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1491] = heapMem[localMem[1456]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3320;
      end

       3320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1491]*6 + localMem[1490]] = localMem[1457];
              updateArrayLength(1, localMem[1491], localMem[1490]);
              ip = 3321;
      end

       3321 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3461;
      end

       3322 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3345;
      end

       3323 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3324;
      end

       3324 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 3325;
      end

       3325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1492] = heapMem[localMem[1456]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3326;
      end

       3326 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1493] = 0; k = arraySizes[localMem[1492]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1492] * NArea + i] == localMem[1449]) localMem[1493] = i + 1;
              end
              ip = 3327;
      end

       3327 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1493] = localMem[1493] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3328;
      end

       3328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1494] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3329;
      end

       3329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1495] = heapMem[localMem[1494]*6 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3330;
      end

       3330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1496] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3331;
      end

       3331 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1497] = heapMem[localMem[1496]*6 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3332;
      end

       3332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1498] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3333;
      end

       3333 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1498]] = localMem[1454];
              ip = 3334;
      end

       3334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1499] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3335;
      end

       3335 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1499]] = localMem[1454];
              ip = 3336;
      end

       3336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1500] = heapMem[localMem[1456]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3337;
      end

       3337 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1500] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1493], localMem[1500], arraySizes[localMem[1500]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1493] && i <= arraySizes[localMem[1500]]) begin
                  heapMem[NArea * localMem[1500] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1500] + localMem[1493]] = localMem[1495];                                    // Insert new value
              arraySizes[localMem[1500]] = arraySizes[localMem[1500]] + 1;                              // Increase array size
              ip = 3338;
      end

       3338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1501] = heapMem[localMem[1456]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3339;
      end

       3339 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1501] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1493], localMem[1501], arraySizes[localMem[1501]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1493] && i <= arraySizes[localMem[1501]]) begin
                  heapMem[NArea * localMem[1501] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1501] + localMem[1493]] = localMem[1497];                                    // Insert new value
              arraySizes[localMem[1501]] = arraySizes[localMem[1501]] + 1;                              // Increase array size
              ip = 3340;
      end

       3340 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1502] = heapMem[localMem[1456]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3341;
      end

       3341 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1503] = localMem[1493] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3342;
      end

       3342 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1502] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1503], localMem[1502], arraySizes[localMem[1502]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1503] && i <= arraySizes[localMem[1502]]) begin
                  heapMem[NArea * localMem[1502] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1502] + localMem[1503]] = localMem[1457];                                    // Insert new value
              arraySizes[localMem[1502]] = arraySizes[localMem[1502]] + 1;                              // Increase array size
              ip = 3343;
      end

       3343 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1456]*6 + 0] = heapMem[localMem[1456]*6 + 0] + 1;
              updateArrayLength(1, localMem[1456], 0);
              ip = 3344;
      end

       3344 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3461;
      end

       3345 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3346;
      end

       3346 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3347;
      end

       3347 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1504] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1504] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1504]] = 0;
              ip = 3348;
      end

       3348 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 0] = localMem[1454];
              updateArrayLength(1, localMem[1504], 0);
              ip = 3349;
      end

       3349 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 2] = 0;
              updateArrayLength(1, localMem[1504], 2);
              ip = 3350;
      end

       3350 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1505] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1505] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1505]] = 0;
              ip = 3351;
      end

       3351 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 4] = localMem[1505];
              updateArrayLength(1, localMem[1504], 4);
              ip = 3352;
      end

       3352 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1506] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1506] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1506]] = 0;
              ip = 3353;
      end

       3353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 5] = localMem[1506];
              updateArrayLength(1, localMem[1504], 5);
              ip = 3354;
      end

       3354 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 6] = 0;
              updateArrayLength(1, localMem[1504], 6);
              ip = 3355;
      end

       3355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 3] = localMem[1452];
              updateArrayLength(1, localMem[1504], 3);
              ip = 3356;
      end

       3356 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1452]*6 + 1] = heapMem[localMem[1452]*6 + 1] + 1;
              updateArrayLength(1, localMem[1452], 1);
              ip = 3357;
      end

       3357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 1] = heapMem[localMem[1452]*6 + 1];
              updateArrayLength(1, localMem[1504], 1);
              ip = 3358;
      end

       3358 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1507] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1507] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1507]] = 0;
              ip = 3359;
      end

       3359 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 0] = localMem[1454];
              updateArrayLength(1, localMem[1507], 0);
              ip = 3360;
      end

       3360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 2] = 0;
              updateArrayLength(1, localMem[1507], 2);
              ip = 3361;
      end

       3361 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1508] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1508] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1508]] = 0;
              ip = 3362;
      end

       3362 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 4] = localMem[1508];
              updateArrayLength(1, localMem[1507], 4);
              ip = 3363;
      end

       3363 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1509] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1509] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1509]] = 0;
              ip = 3364;
      end

       3364 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 5] = localMem[1509];
              updateArrayLength(1, localMem[1507], 5);
              ip = 3365;
      end

       3365 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 6] = 0;
              updateArrayLength(1, localMem[1507], 6);
              ip = 3366;
      end

       3366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 3] = localMem[1452];
              updateArrayLength(1, localMem[1507], 3);
              ip = 3367;
      end

       3367 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1452]*6 + 1] = heapMem[localMem[1452]*6 + 1] + 1;
              updateArrayLength(1, localMem[1452], 1);
              ip = 3368;
      end

       3368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 1] = heapMem[localMem[1452]*6 + 1];
              updateArrayLength(1, localMem[1507], 1);
              ip = 3369;
      end

       3369 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1510] = !heapMem[localMem[1449]*6 + 6];
              ip = 3370;
      end

       3370 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1510] != 0 ? 3422 : 3371;
      end

       3371 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1511] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1511] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1511]] = 0;
              ip = 3372;
      end

       3372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 6] = localMem[1511];
              updateArrayLength(1, localMem[1504], 6);
              ip = 3373;
      end

       3373 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1512] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1512] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1512]] = 0;
              ip = 3374;
      end

       3374 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 6] = localMem[1512];
              updateArrayLength(1, localMem[1507], 6);
              ip = 3375;
      end

       3375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1513] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3376;
      end

       3376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1514] = heapMem[localMem[1504]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3377;
      end

       3377 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1514] + 0 + i] = heapMem[NArea * localMem[1513] + 0 + i];
                  updateArrayLength(1, localMem[1514], 0 + i);
                end
              end
              ip = 3378;
      end

       3378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1515] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3379;
      end

       3379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1516] = heapMem[localMem[1504]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3380;
      end

       3380 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1516] + 0 + i] = heapMem[NArea * localMem[1515] + 0 + i];
                  updateArrayLength(1, localMem[1516], 0 + i);
                end
              end
              ip = 3381;
      end

       3381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1517] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3382;
      end

       3382 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1518] = heapMem[localMem[1504]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3383;
      end

       3383 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1519] = localMem[1454] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3384;
      end

       3384 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1519]) begin
                  heapMem[NArea * localMem[1518] + 0 + i] = heapMem[NArea * localMem[1517] + 0 + i];
                  updateArrayLength(1, localMem[1518], 0 + i);
                end
              end
              ip = 3385;
      end

       3385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1520] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3386;
      end

       3386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1521] = heapMem[localMem[1507]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3387;
      end

       3387 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1521] + 0 + i] = heapMem[NArea * localMem[1520] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1521], 0 + i);
                end
              end
              ip = 3388;
      end

       3388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1522] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3389;
      end

       3389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1523] = heapMem[localMem[1507]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3390;
      end

       3390 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1523] + 0 + i] = heapMem[NArea * localMem[1522] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1523], 0 + i);
                end
              end
              ip = 3391;
      end

       3391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1524] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3392;
      end

       3392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1525] = heapMem[localMem[1507]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3393;
      end

       3393 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1526] = localMem[1454] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3394;
      end

       3394 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1526]) begin
                  heapMem[NArea * localMem[1525] + 0 + i] = heapMem[NArea * localMem[1524] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1525], 0 + i);
                end
              end
              ip = 3395;
      end

       3395 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1527] = heapMem[localMem[1504]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3396;
      end

       3396 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1528] = localMem[1527] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3397;
      end

       3397 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1529] = heapMem[localMem[1504]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3398;
      end

       3398 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3399;
      end

       3399 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1530] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3400;
      end

       3400 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3401;
      end

       3401 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1530] >= localMem[1528] ? 3407 : 3402;
      end

       3402 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1531] = heapMem[localMem[1529]*6 + localMem[1530]];
              updateArrayLength(2, 0, 0);
              ip = 3403;
      end

       3403 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1531]*6 + 2] = localMem[1504];
              updateArrayLength(1, localMem[1531], 2);
              ip = 3404;
      end

       3404 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3405;
      end

       3405 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1530] = localMem[1530] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3406;
      end

       3406 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3400;
      end

       3407 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3408;
      end

       3408 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1532] = heapMem[localMem[1507]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3409;
      end

       3409 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1533] = localMem[1532] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3410;
      end

       3410 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1534] = heapMem[localMem[1507]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3411;
      end

       3411 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3412;
      end

       3412 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1535] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3413;
      end

       3413 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3414;
      end

       3414 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1535] >= localMem[1533] ? 3420 : 3415;
      end

       3415 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1536] = heapMem[localMem[1534]*6 + localMem[1535]];
              updateArrayLength(2, 0, 0);
              ip = 3416;
      end

       3416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1536]*6 + 2] = localMem[1507];
              updateArrayLength(1, localMem[1536], 2);
              ip = 3417;
      end

       3417 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3418;
      end

       3418 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1535] = localMem[1535] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3419;
      end

       3419 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3413;
      end

       3420 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3421;
      end

       3421 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3437;
      end

       3422 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3423;
      end

       3423 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1537] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1537] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1537]] = 0;
              ip = 3424;
      end

       3424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1449]*6 + 6] = localMem[1537];
              updateArrayLength(1, localMem[1449], 6);
              ip = 3425;
      end

       3425 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1538] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3426;
      end

       3426 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1539] = heapMem[localMem[1504]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3427;
      end

       3427 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1539] + 0 + i] = heapMem[NArea * localMem[1538] + 0 + i];
                  updateArrayLength(1, localMem[1539], 0 + i);
                end
              end
              ip = 3428;
      end

       3428 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1540] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3429;
      end

       3429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1541] = heapMem[localMem[1504]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3430;
      end

       3430 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1541] + 0 + i] = heapMem[NArea * localMem[1540] + 0 + i];
                  updateArrayLength(1, localMem[1541], 0 + i);
                end
              end
              ip = 3431;
      end

       3431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1542] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3432;
      end

       3432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1543] = heapMem[localMem[1507]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3433;
      end

       3433 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1543] + 0 + i] = heapMem[NArea * localMem[1542] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1543], 0 + i);
                end
              end
              ip = 3434;
      end

       3434 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1544] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3435;
      end

       3435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1545] = heapMem[localMem[1507]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3436;
      end

       3436 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1545] + 0 + i] = heapMem[NArea * localMem[1544] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1545], 0 + i);
                end
              end
              ip = 3437;
      end

       3437 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3438;
      end

       3438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*6 + 2] = localMem[1449];
              updateArrayLength(1, localMem[1504], 2);
              ip = 3439;
      end

       3439 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*6 + 2] = localMem[1449];
              updateArrayLength(1, localMem[1507], 2);
              ip = 3440;
      end

       3440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1546] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3441;
      end

       3441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1547] = heapMem[localMem[1546]*6 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3442;
      end

       3442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1548] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3443;
      end

       3443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1549] = heapMem[localMem[1548]*6 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3444;
      end

       3444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1550] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3445;
      end

       3445 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1550]*6 + 0] = localMem[1547];
              updateArrayLength(1, localMem[1550], 0);
              ip = 3446;
      end

       3446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1551] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3447;
      end

       3447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1551]*6 + 0] = localMem[1549];
              updateArrayLength(1, localMem[1551], 0);
              ip = 3448;
      end

       3448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1552] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3449;
      end

       3449 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1552]*6 + 0] = localMem[1504];
              updateArrayLength(1, localMem[1552], 0);
              ip = 3450;
      end

       3450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1553] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3451;
      end

       3451 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1553]*6 + 1] = localMem[1507];
              updateArrayLength(1, localMem[1553], 1);
              ip = 3452;
      end

       3452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1449]*6 + 0] = 1;
              updateArrayLength(1, localMem[1449], 0);
              ip = 3453;
      end

       3453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1554] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3454;
      end

       3454 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1554]] = 1;
              ip = 3455;
      end

       3455 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1555] = heapMem[localMem[1449]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3456;
      end

       3456 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1555]] = 1;
              ip = 3457;
      end

       3457 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1556] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3458;
      end

       3458 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1556]] = 2;
              ip = 3459;
      end

       3459 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3461;
      end

       3460 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3466;
      end

       3461 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3462;
      end

       3462 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1450] = 1;
              updateArrayLength(2, 0, 0);
              ip = 3463;
      end

       3463 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3466;
      end

       3464 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3465;
      end

       3465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1450] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3466;
      end

       3466 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3467;
      end

       3467 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3468;
      end

       3468 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3469;
      end

       3469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1557] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3470;
      end

       3470 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3471;
      end

       3471 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1557] >= 99 ? 3969 : 3472;
      end

       3472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1558] = heapMem[localMem[1449]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3473;
      end

       3473 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1559] = localMem[1558] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3474;
      end

       3474 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1560] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3475;
      end

       3475 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1561] = heapMem[localMem[1560]*6 + localMem[1559]];
              updateArrayLength(2, 0, 0);
              ip = 3476;
      end

       3476 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 4 <= localMem[1561] ? 3717 : 3477;
      end

       3477 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1562] = !heapMem[localMem[1449]*6 + 6];
              ip = 3478;
      end

       3478 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1562] == 0 ? 3483 : 3479;
      end

       3479 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 0] = localMem[1449];
              updateArrayLength(1, localMem[1426], 0);
              ip = 3480;
      end

       3480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 1] = 2;
              updateArrayLength(1, localMem[1426], 1);
              ip = 3481;
      end

       3481 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1426]*6 + 2] = localMem[1558] - 1;
              updateArrayLength(1, localMem[1426], 2);
              ip = 3482;
      end

       3482 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3973;
      end

       3483 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3484;
      end

       3484 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1563] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3485;
      end

       3485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1564] = heapMem[localMem[1563]*6 + localMem[1558]];
              updateArrayLength(2, 0, 0);
              ip = 3486;
      end

       3486 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3487;
      end

       3487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1566] = heapMem[localMem[1564]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3488;
      end

       3488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1567] = heapMem[localMem[1564]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3489;
      end

       3489 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1568] = heapMem[localMem[1567]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3490;
      end

       3490 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1566] <  localMem[1568] ? 3710 : 3491;
      end

       3491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1569] = localMem[1568];
              updateArrayLength(2, 0, 0);
              ip = 3492;
      end

       3492 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1569] = localMem[1569] >> 1;
              ip = 3493;
      end

       3493 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1570] = localMem[1569] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3494;
      end

       3494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1571] = heapMem[localMem[1564]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3495;
      end

       3495 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1571] == 0 ? 3592 : 3496;
      end

       3496 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1572] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1572] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1572]] = 0;
              ip = 3497;
      end

       3497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 0] = localMem[1569];
              updateArrayLength(1, localMem[1572], 0);
              ip = 3498;
      end

       3498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 2] = 0;
              updateArrayLength(1, localMem[1572], 2);
              ip = 3499;
      end

       3499 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1573] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1573] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1573]] = 0;
              ip = 3500;
      end

       3500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 4] = localMem[1573];
              updateArrayLength(1, localMem[1572], 4);
              ip = 3501;
      end

       3501 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1574] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1574] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1574]] = 0;
              ip = 3502;
      end

       3502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 5] = localMem[1574];
              updateArrayLength(1, localMem[1572], 5);
              ip = 3503;
      end

       3503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 6] = 0;
              updateArrayLength(1, localMem[1572], 6);
              ip = 3504;
      end

       3504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 3] = localMem[1567];
              updateArrayLength(1, localMem[1572], 3);
              ip = 3505;
      end

       3505 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1567]*6 + 1] = heapMem[localMem[1567]*6 + 1] + 1;
              updateArrayLength(1, localMem[1567], 1);
              ip = 3506;
      end

       3506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 1] = heapMem[localMem[1567]*6 + 1];
              updateArrayLength(1, localMem[1572], 1);
              ip = 3507;
      end

       3507 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1575] = !heapMem[localMem[1564]*6 + 6];
              ip = 3508;
      end

       3508 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1575] != 0 ? 3537 : 3509;
      end

       3509 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1576] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1576] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1576]] = 0;
              ip = 3510;
      end

       3510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 6] = localMem[1576];
              updateArrayLength(1, localMem[1572], 6);
              ip = 3511;
      end

       3511 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1577] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3512;
      end

       3512 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1578] = heapMem[localMem[1572]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3513;
      end

       3513 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1578] + 0 + i] = heapMem[NArea * localMem[1577] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1578], 0 + i);
                end
              end
              ip = 3514;
      end

       3514 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1579] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3515;
      end

       3515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1580] = heapMem[localMem[1572]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3516;
      end

       3516 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1580] + 0 + i] = heapMem[NArea * localMem[1579] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1580], 0 + i);
                end
              end
              ip = 3517;
      end

       3517 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1581] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3518;
      end

       3518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1582] = heapMem[localMem[1572]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3519;
      end

       3519 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1583] = localMem[1569] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3520;
      end

       3520 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1583]) begin
                  heapMem[NArea * localMem[1582] + 0 + i] = heapMem[NArea * localMem[1581] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1582], 0 + i);
                end
              end
              ip = 3521;
      end

       3521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1584] = heapMem[localMem[1572]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3522;
      end

       3522 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1585] = localMem[1584] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3523;
      end

       3523 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1586] = heapMem[localMem[1572]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3524;
      end

       3524 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3525;
      end

       3525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1587] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3526;
      end

       3526 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3527;
      end

       3527 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1587] >= localMem[1585] ? 3533 : 3528;
      end

       3528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1588] = heapMem[localMem[1586]*6 + localMem[1587]];
              updateArrayLength(2, 0, 0);
              ip = 3529;
      end

       3529 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1588]*6 + 2] = localMem[1572];
              updateArrayLength(1, localMem[1588], 2);
              ip = 3530;
      end

       3530 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3531;
      end

       3531 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1587] = localMem[1587] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3532;
      end

       3532 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3526;
      end

       3533 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3534;
      end

       3534 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1589] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3535;
      end

       3535 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1589]] = localMem[1570];
              ip = 3536;
      end

       3536 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3544;
      end

       3537 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3538;
      end

       3538 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1590] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3539;
      end

       3539 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1591] = heapMem[localMem[1572]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3540;
      end

       3540 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1591] + 0 + i] = heapMem[NArea * localMem[1590] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1591], 0 + i);
                end
              end
              ip = 3541;
      end

       3541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1592] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3542;
      end

       3542 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1593] = heapMem[localMem[1572]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3543;
      end

       3543 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1593] + 0 + i] = heapMem[NArea * localMem[1592] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1593], 0 + i);
                end
              end
              ip = 3544;
      end

       3544 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3545;
      end

       3545 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1564]*6 + 0] = localMem[1569];
              updateArrayLength(1, localMem[1564], 0);
              ip = 3546;
      end

       3546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1572]*6 + 2] = localMem[1571];
              updateArrayLength(1, localMem[1572], 2);
              ip = 3547;
      end

       3547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1594] = heapMem[localMem[1571]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3548;
      end

       3548 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1595] = heapMem[localMem[1571]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3549;
      end

       3549 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1596] = heapMem[localMem[1595]*6 + localMem[1594]];
              updateArrayLength(2, 0, 0);
              ip = 3550;
      end

       3550 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1596] != localMem[1564] ? 3569 : 3551;
      end

       3551 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1597] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3552;
      end

       3552 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1598] = heapMem[localMem[1597]*6 + localMem[1569]];
              updateArrayLength(2, 0, 0);
              ip = 3553;
      end

       3553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1599] = heapMem[localMem[1571]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3554;
      end

       3554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1599]*6 + localMem[1594]] = localMem[1598];
              updateArrayLength(1, localMem[1599], localMem[1594]);
              ip = 3555;
      end

       3555 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1600] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3556;
      end

       3556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1601] = heapMem[localMem[1600]*6 + localMem[1569]];
              updateArrayLength(2, 0, 0);
              ip = 3557;
      end

       3557 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1602] = heapMem[localMem[1571]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3558;
      end

       3558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1602]*6 + localMem[1594]] = localMem[1601];
              updateArrayLength(1, localMem[1602], localMem[1594]);
              ip = 3559;
      end

       3559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1603] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3560;
      end

       3560 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1603]] = localMem[1569];
              ip = 3561;
      end

       3561 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1604] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3562;
      end

       3562 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1604]] = localMem[1569];
              ip = 3563;
      end

       3563 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1605] = localMem[1594] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3564;
      end

       3564 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1571]*6 + 0] = localMem[1605];
              updateArrayLength(1, localMem[1571], 0);
              ip = 3565;
      end

       3565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1606] = heapMem[localMem[1571]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3566;
      end

       3566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1606]*6 + localMem[1605]] = localMem[1572];
              updateArrayLength(1, localMem[1606], localMem[1605]);
              ip = 3567;
      end

       3567 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3707;
      end

       3568 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3591;
      end

       3569 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3570;
      end

       3570 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 3571;
      end

       3571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1607] = heapMem[localMem[1571]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3572;
      end

       3572 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1608] = 0; k = arraySizes[localMem[1607]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1607] * NArea + i] == localMem[1564]) localMem[1608] = i + 1;
              end
              ip = 3573;
      end

       3573 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1608] = localMem[1608] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3574;
      end

       3574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1609] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3575;
      end

       3575 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1610] = heapMem[localMem[1609]*6 + localMem[1569]];
              updateArrayLength(2, 0, 0);
              ip = 3576;
      end

       3576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1611] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3577;
      end

       3577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1612] = heapMem[localMem[1611]*6 + localMem[1569]];
              updateArrayLength(2, 0, 0);
              ip = 3578;
      end

       3578 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1613] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3579;
      end

       3579 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1613]] = localMem[1569];
              ip = 3580;
      end

       3580 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1614] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3581;
      end

       3581 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1614]] = localMem[1569];
              ip = 3582;
      end

       3582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1615] = heapMem[localMem[1571]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3583;
      end

       3583 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1615] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1608], localMem[1615], arraySizes[localMem[1615]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1608] && i <= arraySizes[localMem[1615]]) begin
                  heapMem[NArea * localMem[1615] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1615] + localMem[1608]] = localMem[1610];                                    // Insert new value
              arraySizes[localMem[1615]] = arraySizes[localMem[1615]] + 1;                              // Increase array size
              ip = 3584;
      end

       3584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1616] = heapMem[localMem[1571]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3585;
      end

       3585 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1616] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1608], localMem[1616], arraySizes[localMem[1616]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1608] && i <= arraySizes[localMem[1616]]) begin
                  heapMem[NArea * localMem[1616] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1616] + localMem[1608]] = localMem[1612];                                    // Insert new value
              arraySizes[localMem[1616]] = arraySizes[localMem[1616]] + 1;                              // Increase array size
              ip = 3586;
      end

       3586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1617] = heapMem[localMem[1571]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3587;
      end

       3587 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1618] = localMem[1608] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3588;
      end

       3588 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1617] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1618], localMem[1617], arraySizes[localMem[1617]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1618] && i <= arraySizes[localMem[1617]]) begin
                  heapMem[NArea * localMem[1617] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1617] + localMem[1618]] = localMem[1572];                                    // Insert new value
              arraySizes[localMem[1617]] = arraySizes[localMem[1617]] + 1;                              // Increase array size
              ip = 3589;
      end

       3589 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1571]*6 + 0] = heapMem[localMem[1571]*6 + 0] + 1;
              updateArrayLength(1, localMem[1571], 0);
              ip = 3590;
      end

       3590 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3707;
      end

       3591 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3592;
      end

       3592 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3593;
      end

       3593 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1619] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1619] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1619]] = 0;
              ip = 3594;
      end

       3594 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 0] = localMem[1569];
              updateArrayLength(1, localMem[1619], 0);
              ip = 3595;
      end

       3595 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 2] = 0;
              updateArrayLength(1, localMem[1619], 2);
              ip = 3596;
      end

       3596 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1620] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1620] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1620]] = 0;
              ip = 3597;
      end

       3597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 4] = localMem[1620];
              updateArrayLength(1, localMem[1619], 4);
              ip = 3598;
      end

       3598 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1621] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1621] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1621]] = 0;
              ip = 3599;
      end

       3599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 5] = localMem[1621];
              updateArrayLength(1, localMem[1619], 5);
              ip = 3600;
      end

       3600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 6] = 0;
              updateArrayLength(1, localMem[1619], 6);
              ip = 3601;
      end

       3601 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 3] = localMem[1567];
              updateArrayLength(1, localMem[1619], 3);
              ip = 3602;
      end

       3602 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1567]*6 + 1] = heapMem[localMem[1567]*6 + 1] + 1;
              updateArrayLength(1, localMem[1567], 1);
              ip = 3603;
      end

       3603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 1] = heapMem[localMem[1567]*6 + 1];
              updateArrayLength(1, localMem[1619], 1);
              ip = 3604;
      end

       3604 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1622] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1622] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1622]] = 0;
              ip = 3605;
      end

       3605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 0] = localMem[1569];
              updateArrayLength(1, localMem[1622], 0);
              ip = 3606;
      end

       3606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 2] = 0;
              updateArrayLength(1, localMem[1622], 2);
              ip = 3607;
      end

       3607 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1623] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1623] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1623]] = 0;
              ip = 3608;
      end

       3608 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 4] = localMem[1623];
              updateArrayLength(1, localMem[1622], 4);
              ip = 3609;
      end

       3609 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1624] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1624] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1624]] = 0;
              ip = 3610;
      end

       3610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 5] = localMem[1624];
              updateArrayLength(1, localMem[1622], 5);
              ip = 3611;
      end

       3611 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 6] = 0;
              updateArrayLength(1, localMem[1622], 6);
              ip = 3612;
      end

       3612 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 3] = localMem[1567];
              updateArrayLength(1, localMem[1622], 3);
              ip = 3613;
      end

       3613 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1567]*6 + 1] = heapMem[localMem[1567]*6 + 1] + 1;
              updateArrayLength(1, localMem[1567], 1);
              ip = 3614;
      end

       3614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 1] = heapMem[localMem[1567]*6 + 1];
              updateArrayLength(1, localMem[1622], 1);
              ip = 3615;
      end

       3615 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1625] = !heapMem[localMem[1564]*6 + 6];
              ip = 3616;
      end

       3616 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1625] != 0 ? 3668 : 3617;
      end

       3617 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1626] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1626] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1626]] = 0;
              ip = 3618;
      end

       3618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 6] = localMem[1626];
              updateArrayLength(1, localMem[1619], 6);
              ip = 3619;
      end

       3619 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1627] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1627] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1627]] = 0;
              ip = 3620;
      end

       3620 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 6] = localMem[1627];
              updateArrayLength(1, localMem[1622], 6);
              ip = 3621;
      end

       3621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1628] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3622;
      end

       3622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1629] = heapMem[localMem[1619]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3623;
      end

       3623 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1629] + 0 + i] = heapMem[NArea * localMem[1628] + 0 + i];
                  updateArrayLength(1, localMem[1629], 0 + i);
                end
              end
              ip = 3624;
      end

       3624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1630] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3625;
      end

       3625 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1631] = heapMem[localMem[1619]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3626;
      end

       3626 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1631] + 0 + i] = heapMem[NArea * localMem[1630] + 0 + i];
                  updateArrayLength(1, localMem[1631], 0 + i);
                end
              end
              ip = 3627;
      end

       3627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1632] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3628;
      end

       3628 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1633] = heapMem[localMem[1619]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3629;
      end

       3629 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1634] = localMem[1569] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3630;
      end

       3630 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1634]) begin
                  heapMem[NArea * localMem[1633] + 0 + i] = heapMem[NArea * localMem[1632] + 0 + i];
                  updateArrayLength(1, localMem[1633], 0 + i);
                end
              end
              ip = 3631;
      end

       3631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1635] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3632;
      end

       3632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1636] = heapMem[localMem[1622]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3633;
      end

       3633 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1636] + 0 + i] = heapMem[NArea * localMem[1635] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1636], 0 + i);
                end
              end
              ip = 3634;
      end

       3634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1637] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3635;
      end

       3635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1638] = heapMem[localMem[1622]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3636;
      end

       3636 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1638] + 0 + i] = heapMem[NArea * localMem[1637] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1638], 0 + i);
                end
              end
              ip = 3637;
      end

       3637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1639] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3638;
      end

       3638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1640] = heapMem[localMem[1622]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3639;
      end

       3639 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1641] = localMem[1569] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3640;
      end

       3640 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1641]) begin
                  heapMem[NArea * localMem[1640] + 0 + i] = heapMem[NArea * localMem[1639] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1640], 0 + i);
                end
              end
              ip = 3641;
      end

       3641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1642] = heapMem[localMem[1619]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3642;
      end

       3642 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1643] = localMem[1642] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3643;
      end

       3643 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1644] = heapMem[localMem[1619]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3644;
      end

       3644 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3645;
      end

       3645 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1645] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3646;
      end

       3646 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3647;
      end

       3647 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1645] >= localMem[1643] ? 3653 : 3648;
      end

       3648 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1646] = heapMem[localMem[1644]*6 + localMem[1645]];
              updateArrayLength(2, 0, 0);
              ip = 3649;
      end

       3649 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1646]*6 + 2] = localMem[1619];
              updateArrayLength(1, localMem[1646], 2);
              ip = 3650;
      end

       3650 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3651;
      end

       3651 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1645] = localMem[1645] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3652;
      end

       3652 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3646;
      end

       3653 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3654;
      end

       3654 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1647] = heapMem[localMem[1622]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3655;
      end

       3655 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1648] = localMem[1647] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3656;
      end

       3656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1649] = heapMem[localMem[1622]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3657;
      end

       3657 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3658;
      end

       3658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1650] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3659;
      end

       3659 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3660;
      end

       3660 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1650] >= localMem[1648] ? 3666 : 3661;
      end

       3661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1651] = heapMem[localMem[1649]*6 + localMem[1650]];
              updateArrayLength(2, 0, 0);
              ip = 3662;
      end

       3662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1651]*6 + 2] = localMem[1622];
              updateArrayLength(1, localMem[1651], 2);
              ip = 3663;
      end

       3663 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3664;
      end

       3664 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1650] = localMem[1650] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3665;
      end

       3665 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3659;
      end

       3666 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3667;
      end

       3667 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3683;
      end

       3668 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3669;
      end

       3669 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1652] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1652] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1652]] = 0;
              ip = 3670;
      end

       3670 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1564]*6 + 6] = localMem[1652];
              updateArrayLength(1, localMem[1564], 6);
              ip = 3671;
      end

       3671 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1653] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3672;
      end

       3672 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1654] = heapMem[localMem[1619]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3673;
      end

       3673 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1654] + 0 + i] = heapMem[NArea * localMem[1653] + 0 + i];
                  updateArrayLength(1, localMem[1654], 0 + i);
                end
              end
              ip = 3674;
      end

       3674 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1655] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3675;
      end

       3675 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1656] = heapMem[localMem[1619]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3676;
      end

       3676 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1656] + 0 + i] = heapMem[NArea * localMem[1655] + 0 + i];
                  updateArrayLength(1, localMem[1656], 0 + i);
                end
              end
              ip = 3677;
      end

       3677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1657] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3678;
      end

       3678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1658] = heapMem[localMem[1622]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3679;
      end

       3679 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1658] + 0 + i] = heapMem[NArea * localMem[1657] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1658], 0 + i);
                end
              end
              ip = 3680;
      end

       3680 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1659] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3681;
      end

       3681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1660] = heapMem[localMem[1622]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3682;
      end

       3682 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1569]) begin
                  heapMem[NArea * localMem[1660] + 0 + i] = heapMem[NArea * localMem[1659] + localMem[1570] + i];
                  updateArrayLength(1, localMem[1660], 0 + i);
                end
              end
              ip = 3683;
      end

       3683 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3684;
      end

       3684 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1619]*6 + 2] = localMem[1564];
              updateArrayLength(1, localMem[1619], 2);
              ip = 3685;
      end

       3685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1622]*6 + 2] = localMem[1564];
              updateArrayLength(1, localMem[1622], 2);
              ip = 3686;
      end

       3686 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1661] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3687;
      end

       3687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1662] = heapMem[localMem[1661]*6 + localMem[1569]];
              updateArrayLength(2, 0, 0);
              ip = 3688;
      end

       3688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1663] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3689;
      end

       3689 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1664] = heapMem[localMem[1663]*6 + localMem[1569]];
              updateArrayLength(2, 0, 0);
              ip = 3690;
      end

       3690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1665] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3691;
      end

       3691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1665]*6 + 0] = localMem[1662];
              updateArrayLength(1, localMem[1665], 0);
              ip = 3692;
      end

       3692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1666] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3693;
      end

       3693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1666]*6 + 0] = localMem[1664];
              updateArrayLength(1, localMem[1666], 0);
              ip = 3694;
      end

       3694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1667] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3695;
      end

       3695 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1667]*6 + 0] = localMem[1619];
              updateArrayLength(1, localMem[1667], 0);
              ip = 3696;
      end

       3696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1668] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3697;
      end

       3697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1668]*6 + 1] = localMem[1622];
              updateArrayLength(1, localMem[1668], 1);
              ip = 3698;
      end

       3698 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1564]*6 + 0] = 1;
              updateArrayLength(1, localMem[1564], 0);
              ip = 3699;
      end

       3699 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1669] = heapMem[localMem[1564]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3700;
      end

       3700 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1669]] = 1;
              ip = 3701;
      end

       3701 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1670] = heapMem[localMem[1564]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3702;
      end

       3702 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1670]] = 1;
              ip = 3703;
      end

       3703 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1671] = heapMem[localMem[1564]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3704;
      end

       3704 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1671]] = 2;
              ip = 3705;
      end

       3705 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3707;
      end

       3706 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3712;
      end

       3707 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3708;
      end

       3708 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1565] = 1;
              updateArrayLength(2, 0, 0);
              ip = 3709;
      end

       3709 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3712;
      end

       3710 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3711;
      end

       3711 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1565] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3712;
      end

       3712 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3713;
      end

       3713 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1565] != 0 ? 3715 : 3714;
      end

       3714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1449] = localMem[1564];
              updateArrayLength(2, 0, 0);
              ip = 3715;
      end

       3715 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3716;
      end

       3716 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3966;
      end

       3717 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3718;
      end

       3718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1672] = heapMem[localMem[1449]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3719;
      end

       3719 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1673] = 0; k = arraySizes[localMem[1672]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1672] * NArea + i] == 4) localMem[1673] = i + 1;
              end
              ip = 3720;
      end

       3720 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1673] == 0 ? 3725 : 3721;
      end

       3721 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 0] = localMem[1449];
              updateArrayLength(1, localMem[1426], 0);
              ip = 3722;
      end

       3722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 1] = 1;
              updateArrayLength(1, localMem[1426], 1);
              ip = 3723;
      end

       3723 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1426]*6 + 2] = localMem[1673] - 1;
              updateArrayLength(1, localMem[1426], 2);
              ip = 3724;
      end

       3724 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3973;
      end

       3725 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3726;
      end

       3726 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[1672]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1672] * NArea + i] < 4) j = j + 1;
              end
              localMem[1674] = j;
              ip = 3727;
      end

       3727 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1675] = !heapMem[localMem[1449]*6 + 6];
              ip = 3728;
      end

       3728 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1675] == 0 ? 3733 : 3729;
      end

       3729 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 0] = localMem[1449];
              updateArrayLength(1, localMem[1426], 0);
              ip = 3730;
      end

       3730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 1] = 0;
              updateArrayLength(1, localMem[1426], 1);
              ip = 3731;
      end

       3731 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*6 + 2] = localMem[1674];
              updateArrayLength(1, localMem[1426], 2);
              ip = 3732;
      end

       3732 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3973;
      end

       3733 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3734;
      end

       3734 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1676] = heapMem[localMem[1449]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3735;
      end

       3735 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1677] = heapMem[localMem[1676]*6 + localMem[1674]];
              updateArrayLength(2, 0, 0);
              ip = 3736;
      end

       3736 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3737;
      end

       3737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1679] = heapMem[localMem[1677]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3738;
      end

       3738 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1680] = heapMem[localMem[1677]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3739;
      end

       3739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1681] = heapMem[localMem[1680]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3740;
      end

       3740 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1679] <  localMem[1681] ? 3960 : 3741;
      end

       3741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1682] = localMem[1681];
              updateArrayLength(2, 0, 0);
              ip = 3742;
      end

       3742 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1682] = localMem[1682] >> 1;
              ip = 3743;
      end

       3743 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1683] = localMem[1682] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3744;
      end

       3744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1684] = heapMem[localMem[1677]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3745;
      end

       3745 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1684] == 0 ? 3842 : 3746;
      end

       3746 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1685] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1685] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1685]] = 0;
              ip = 3747;
      end

       3747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 0] = localMem[1682];
              updateArrayLength(1, localMem[1685], 0);
              ip = 3748;
      end

       3748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 2] = 0;
              updateArrayLength(1, localMem[1685], 2);
              ip = 3749;
      end

       3749 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1686] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1686] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1686]] = 0;
              ip = 3750;
      end

       3750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 4] = localMem[1686];
              updateArrayLength(1, localMem[1685], 4);
              ip = 3751;
      end

       3751 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1687] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1687] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1687]] = 0;
              ip = 3752;
      end

       3752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 5] = localMem[1687];
              updateArrayLength(1, localMem[1685], 5);
              ip = 3753;
      end

       3753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 6] = 0;
              updateArrayLength(1, localMem[1685], 6);
              ip = 3754;
      end

       3754 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 3] = localMem[1680];
              updateArrayLength(1, localMem[1685], 3);
              ip = 3755;
      end

       3755 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1680]*6 + 1] = heapMem[localMem[1680]*6 + 1] + 1;
              updateArrayLength(1, localMem[1680], 1);
              ip = 3756;
      end

       3756 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 1] = heapMem[localMem[1680]*6 + 1];
              updateArrayLength(1, localMem[1685], 1);
              ip = 3757;
      end

       3757 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1688] = !heapMem[localMem[1677]*6 + 6];
              ip = 3758;
      end

       3758 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1688] != 0 ? 3787 : 3759;
      end

       3759 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1689] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1689] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1689]] = 0;
              ip = 3760;
      end

       3760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 6] = localMem[1689];
              updateArrayLength(1, localMem[1685], 6);
              ip = 3761;
      end

       3761 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1690] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3762;
      end

       3762 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1691] = heapMem[localMem[1685]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3763;
      end

       3763 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1691] + 0 + i] = heapMem[NArea * localMem[1690] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1691], 0 + i);
                end
              end
              ip = 3764;
      end

       3764 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1692] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3765;
      end

       3765 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1693] = heapMem[localMem[1685]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3766;
      end

       3766 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1693] + 0 + i] = heapMem[NArea * localMem[1692] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1693], 0 + i);
                end
              end
              ip = 3767;
      end

       3767 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1694] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3768;
      end

       3768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1695] = heapMem[localMem[1685]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3769;
      end

       3769 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1696] = localMem[1682] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3770;
      end

       3770 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1696]) begin
                  heapMem[NArea * localMem[1695] + 0 + i] = heapMem[NArea * localMem[1694] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1695], 0 + i);
                end
              end
              ip = 3771;
      end

       3771 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1697] = heapMem[localMem[1685]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3772;
      end

       3772 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1698] = localMem[1697] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3773;
      end

       3773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1699] = heapMem[localMem[1685]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3774;
      end

       3774 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3775;
      end

       3775 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1700] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3776;
      end

       3776 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3777;
      end

       3777 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1700] >= localMem[1698] ? 3783 : 3778;
      end

       3778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1701] = heapMem[localMem[1699]*6 + localMem[1700]];
              updateArrayLength(2, 0, 0);
              ip = 3779;
      end

       3779 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1701]*6 + 2] = localMem[1685];
              updateArrayLength(1, localMem[1701], 2);
              ip = 3780;
      end

       3780 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3781;
      end

       3781 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1700] = localMem[1700] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3782;
      end

       3782 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3776;
      end

       3783 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3784;
      end

       3784 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1702] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3785;
      end

       3785 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1702]] = localMem[1683];
              ip = 3786;
      end

       3786 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3794;
      end

       3787 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3788;
      end

       3788 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1703] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3789;
      end

       3789 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1704] = heapMem[localMem[1685]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3790;
      end

       3790 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1704] + 0 + i] = heapMem[NArea * localMem[1703] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1704], 0 + i);
                end
              end
              ip = 3791;
      end

       3791 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1705] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3792;
      end

       3792 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1706] = heapMem[localMem[1685]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3793;
      end

       3793 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1706] + 0 + i] = heapMem[NArea * localMem[1705] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1706], 0 + i);
                end
              end
              ip = 3794;
      end

       3794 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3795;
      end

       3795 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1677]*6 + 0] = localMem[1682];
              updateArrayLength(1, localMem[1677], 0);
              ip = 3796;
      end

       3796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1685]*6 + 2] = localMem[1684];
              updateArrayLength(1, localMem[1685], 2);
              ip = 3797;
      end

       3797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1707] = heapMem[localMem[1684]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3798;
      end

       3798 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1708] = heapMem[localMem[1684]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3799;
      end

       3799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1709] = heapMem[localMem[1708]*6 + localMem[1707]];
              updateArrayLength(2, 0, 0);
              ip = 3800;
      end

       3800 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1709] != localMem[1677] ? 3819 : 3801;
      end

       3801 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1710] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3802;
      end

       3802 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1711] = heapMem[localMem[1710]*6 + localMem[1682]];
              updateArrayLength(2, 0, 0);
              ip = 3803;
      end

       3803 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1712] = heapMem[localMem[1684]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3804;
      end

       3804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1712]*6 + localMem[1707]] = localMem[1711];
              updateArrayLength(1, localMem[1712], localMem[1707]);
              ip = 3805;
      end

       3805 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1713] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3806;
      end

       3806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1714] = heapMem[localMem[1713]*6 + localMem[1682]];
              updateArrayLength(2, 0, 0);
              ip = 3807;
      end

       3807 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1715] = heapMem[localMem[1684]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3808;
      end

       3808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1715]*6 + localMem[1707]] = localMem[1714];
              updateArrayLength(1, localMem[1715], localMem[1707]);
              ip = 3809;
      end

       3809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1716] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3810;
      end

       3810 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1716]] = localMem[1682];
              ip = 3811;
      end

       3811 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1717] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3812;
      end

       3812 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1717]] = localMem[1682];
              ip = 3813;
      end

       3813 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1718] = localMem[1707] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3814;
      end

       3814 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1684]*6 + 0] = localMem[1718];
              updateArrayLength(1, localMem[1684], 0);
              ip = 3815;
      end

       3815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1719] = heapMem[localMem[1684]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3816;
      end

       3816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1719]*6 + localMem[1718]] = localMem[1685];
              updateArrayLength(1, localMem[1719], localMem[1718]);
              ip = 3817;
      end

       3817 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3957;
      end

       3818 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3841;
      end

       3819 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3820;
      end

       3820 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 3821;
      end

       3821 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1720] = heapMem[localMem[1684]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3822;
      end

       3822 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1721] = 0; k = arraySizes[localMem[1720]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1720] * NArea + i] == localMem[1677]) localMem[1721] = i + 1;
              end
              ip = 3823;
      end

       3823 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1721] = localMem[1721] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3824;
      end

       3824 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1722] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3825;
      end

       3825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1723] = heapMem[localMem[1722]*6 + localMem[1682]];
              updateArrayLength(2, 0, 0);
              ip = 3826;
      end

       3826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1724] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3827;
      end

       3827 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1725] = heapMem[localMem[1724]*6 + localMem[1682]];
              updateArrayLength(2, 0, 0);
              ip = 3828;
      end

       3828 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1726] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3829;
      end

       3829 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1726]] = localMem[1682];
              ip = 3830;
      end

       3830 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1727] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3831;
      end

       3831 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1727]] = localMem[1682];
              ip = 3832;
      end

       3832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1728] = heapMem[localMem[1684]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3833;
      end

       3833 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1728] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1721], localMem[1728], arraySizes[localMem[1728]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1721] && i <= arraySizes[localMem[1728]]) begin
                  heapMem[NArea * localMem[1728] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1728] + localMem[1721]] = localMem[1723];                                    // Insert new value
              arraySizes[localMem[1728]] = arraySizes[localMem[1728]] + 1;                              // Increase array size
              ip = 3834;
      end

       3834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1729] = heapMem[localMem[1684]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3835;
      end

       3835 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1729] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1721], localMem[1729], arraySizes[localMem[1729]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1721] && i <= arraySizes[localMem[1729]]) begin
                  heapMem[NArea * localMem[1729] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1729] + localMem[1721]] = localMem[1725];                                    // Insert new value
              arraySizes[localMem[1729]] = arraySizes[localMem[1729]] + 1;                              // Increase array size
              ip = 3836;
      end

       3836 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1730] = heapMem[localMem[1684]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3837;
      end

       3837 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1731] = localMem[1721] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3838;
      end

       3838 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1730] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1731], localMem[1730], arraySizes[localMem[1730]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1731] && i <= arraySizes[localMem[1730]]) begin
                  heapMem[NArea * localMem[1730] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1730] + localMem[1731]] = localMem[1685];                                    // Insert new value
              arraySizes[localMem[1730]] = arraySizes[localMem[1730]] + 1;                              // Increase array size
              ip = 3839;
      end

       3839 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1684]*6 + 0] = heapMem[localMem[1684]*6 + 0] + 1;
              updateArrayLength(1, localMem[1684], 0);
              ip = 3840;
      end

       3840 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3957;
      end

       3841 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3842;
      end

       3842 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3843;
      end

       3843 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1732] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1732] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1732]] = 0;
              ip = 3844;
      end

       3844 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 0] = localMem[1682];
              updateArrayLength(1, localMem[1732], 0);
              ip = 3845;
      end

       3845 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 2] = 0;
              updateArrayLength(1, localMem[1732], 2);
              ip = 3846;
      end

       3846 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1733] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1733] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1733]] = 0;
              ip = 3847;
      end

       3847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 4] = localMem[1733];
              updateArrayLength(1, localMem[1732], 4);
              ip = 3848;
      end

       3848 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1734] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1734] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1734]] = 0;
              ip = 3849;
      end

       3849 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 5] = localMem[1734];
              updateArrayLength(1, localMem[1732], 5);
              ip = 3850;
      end

       3850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 6] = 0;
              updateArrayLength(1, localMem[1732], 6);
              ip = 3851;
      end

       3851 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 3] = localMem[1680];
              updateArrayLength(1, localMem[1732], 3);
              ip = 3852;
      end

       3852 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1680]*6 + 1] = heapMem[localMem[1680]*6 + 1] + 1;
              updateArrayLength(1, localMem[1680], 1);
              ip = 3853;
      end

       3853 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 1] = heapMem[localMem[1680]*6 + 1];
              updateArrayLength(1, localMem[1732], 1);
              ip = 3854;
      end

       3854 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1735] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1735] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1735]] = 0;
              ip = 3855;
      end

       3855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 0] = localMem[1682];
              updateArrayLength(1, localMem[1735], 0);
              ip = 3856;
      end

       3856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 2] = 0;
              updateArrayLength(1, localMem[1735], 2);
              ip = 3857;
      end

       3857 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1736] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1736] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1736]] = 0;
              ip = 3858;
      end

       3858 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 4] = localMem[1736];
              updateArrayLength(1, localMem[1735], 4);
              ip = 3859;
      end

       3859 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1737] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1737] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1737]] = 0;
              ip = 3860;
      end

       3860 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 5] = localMem[1737];
              updateArrayLength(1, localMem[1735], 5);
              ip = 3861;
      end

       3861 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 6] = 0;
              updateArrayLength(1, localMem[1735], 6);
              ip = 3862;
      end

       3862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 3] = localMem[1680];
              updateArrayLength(1, localMem[1735], 3);
              ip = 3863;
      end

       3863 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1680]*6 + 1] = heapMem[localMem[1680]*6 + 1] + 1;
              updateArrayLength(1, localMem[1680], 1);
              ip = 3864;
      end

       3864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 1] = heapMem[localMem[1680]*6 + 1];
              updateArrayLength(1, localMem[1735], 1);
              ip = 3865;
      end

       3865 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1738] = !heapMem[localMem[1677]*6 + 6];
              ip = 3866;
      end

       3866 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1738] != 0 ? 3918 : 3867;
      end

       3867 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1739] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1739] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1739]] = 0;
              ip = 3868;
      end

       3868 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 6] = localMem[1739];
              updateArrayLength(1, localMem[1732], 6);
              ip = 3869;
      end

       3869 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1740] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1740] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1740]] = 0;
              ip = 3870;
      end

       3870 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 6] = localMem[1740];
              updateArrayLength(1, localMem[1735], 6);
              ip = 3871;
      end

       3871 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1741] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3872;
      end

       3872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1742] = heapMem[localMem[1732]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3873;
      end

       3873 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1742] + 0 + i] = heapMem[NArea * localMem[1741] + 0 + i];
                  updateArrayLength(1, localMem[1742], 0 + i);
                end
              end
              ip = 3874;
      end

       3874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1743] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3875;
      end

       3875 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1744] = heapMem[localMem[1732]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3876;
      end

       3876 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1744] + 0 + i] = heapMem[NArea * localMem[1743] + 0 + i];
                  updateArrayLength(1, localMem[1744], 0 + i);
                end
              end
              ip = 3877;
      end

       3877 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1745] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3878;
      end

       3878 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1746] = heapMem[localMem[1732]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3879;
      end

       3879 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1747] = localMem[1682] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3880;
      end

       3880 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1747]) begin
                  heapMem[NArea * localMem[1746] + 0 + i] = heapMem[NArea * localMem[1745] + 0 + i];
                  updateArrayLength(1, localMem[1746], 0 + i);
                end
              end
              ip = 3881;
      end

       3881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1748] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3882;
      end

       3882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1749] = heapMem[localMem[1735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3883;
      end

       3883 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1749] + 0 + i] = heapMem[NArea * localMem[1748] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1749], 0 + i);
                end
              end
              ip = 3884;
      end

       3884 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1750] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3885;
      end

       3885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1751] = heapMem[localMem[1735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3886;
      end

       3886 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1751] + 0 + i] = heapMem[NArea * localMem[1750] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1751], 0 + i);
                end
              end
              ip = 3887;
      end

       3887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1752] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3888;
      end

       3888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1753] = heapMem[localMem[1735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3889;
      end

       3889 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1754] = localMem[1682] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3890;
      end

       3890 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1754]) begin
                  heapMem[NArea * localMem[1753] + 0 + i] = heapMem[NArea * localMem[1752] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1753], 0 + i);
                end
              end
              ip = 3891;
      end

       3891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1755] = heapMem[localMem[1732]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3892;
      end

       3892 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1756] = localMem[1755] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3893;
      end

       3893 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1757] = heapMem[localMem[1732]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3894;
      end

       3894 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3895;
      end

       3895 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1758] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3896;
      end

       3896 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3897;
      end

       3897 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1758] >= localMem[1756] ? 3903 : 3898;
      end

       3898 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1759] = heapMem[localMem[1757]*6 + localMem[1758]];
              updateArrayLength(2, 0, 0);
              ip = 3899;
      end

       3899 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1759]*6 + 2] = localMem[1732];
              updateArrayLength(1, localMem[1759], 2);
              ip = 3900;
      end

       3900 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3901;
      end

       3901 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1758] = localMem[1758] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3902;
      end

       3902 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3896;
      end

       3903 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3904;
      end

       3904 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1760] = heapMem[localMem[1735]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3905;
      end

       3905 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1761] = localMem[1760] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3906;
      end

       3906 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1762] = heapMem[localMem[1735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3907;
      end

       3907 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3908;
      end

       3908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1763] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3909;
      end

       3909 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3910;
      end

       3910 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1763] >= localMem[1761] ? 3916 : 3911;
      end

       3911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1764] = heapMem[localMem[1762]*6 + localMem[1763]];
              updateArrayLength(2, 0, 0);
              ip = 3912;
      end

       3912 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1764]*6 + 2] = localMem[1735];
              updateArrayLength(1, localMem[1764], 2);
              ip = 3913;
      end

       3913 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3914;
      end

       3914 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1763] = localMem[1763] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3915;
      end

       3915 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3909;
      end

       3916 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3917;
      end

       3917 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3933;
      end

       3918 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3919;
      end

       3919 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1765] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1765] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1765]] = 0;
              ip = 3920;
      end

       3920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1677]*6 + 6] = localMem[1765];
              updateArrayLength(1, localMem[1677], 6);
              ip = 3921;
      end

       3921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1766] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3922;
      end

       3922 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1767] = heapMem[localMem[1732]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3923;
      end

       3923 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1767] + 0 + i] = heapMem[NArea * localMem[1766] + 0 + i];
                  updateArrayLength(1, localMem[1767], 0 + i);
                end
              end
              ip = 3924;
      end

       3924 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1768] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3925;
      end

       3925 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1769] = heapMem[localMem[1732]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3926;
      end

       3926 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1769] + 0 + i] = heapMem[NArea * localMem[1768] + 0 + i];
                  updateArrayLength(1, localMem[1769], 0 + i);
                end
              end
              ip = 3927;
      end

       3927 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1770] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3928;
      end

       3928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1771] = heapMem[localMem[1735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3929;
      end

       3929 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1771] + 0 + i] = heapMem[NArea * localMem[1770] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1771], 0 + i);
                end
              end
              ip = 3930;
      end

       3930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1772] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3931;
      end

       3931 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1773] = heapMem[localMem[1735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3932;
      end

       3932 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1682]) begin
                  heapMem[NArea * localMem[1773] + 0 + i] = heapMem[NArea * localMem[1772] + localMem[1683] + i];
                  updateArrayLength(1, localMem[1773], 0 + i);
                end
              end
              ip = 3933;
      end

       3933 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3934;
      end

       3934 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1732]*6 + 2] = localMem[1677];
              updateArrayLength(1, localMem[1732], 2);
              ip = 3935;
      end

       3935 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1735]*6 + 2] = localMem[1677];
              updateArrayLength(1, localMem[1735], 2);
              ip = 3936;
      end

       3936 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1774] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3937;
      end

       3937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1775] = heapMem[localMem[1774]*6 + localMem[1682]];
              updateArrayLength(2, 0, 0);
              ip = 3938;
      end

       3938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1776] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3939;
      end

       3939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1777] = heapMem[localMem[1776]*6 + localMem[1682]];
              updateArrayLength(2, 0, 0);
              ip = 3940;
      end

       3940 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1778] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3941;
      end

       3941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1778]*6 + 0] = localMem[1775];
              updateArrayLength(1, localMem[1778], 0);
              ip = 3942;
      end

       3942 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1779] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3943;
      end

       3943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1779]*6 + 0] = localMem[1777];
              updateArrayLength(1, localMem[1779], 0);
              ip = 3944;
      end

       3944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1780] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3945;
      end

       3945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1780]*6 + 0] = localMem[1732];
              updateArrayLength(1, localMem[1780], 0);
              ip = 3946;
      end

       3946 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1781] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3947;
      end

       3947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1781]*6 + 1] = localMem[1735];
              updateArrayLength(1, localMem[1781], 1);
              ip = 3948;
      end

       3948 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1677]*6 + 0] = 1;
              updateArrayLength(1, localMem[1677], 0);
              ip = 3949;
      end

       3949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1782] = heapMem[localMem[1677]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3950;
      end

       3950 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1782]] = 1;
              ip = 3951;
      end

       3951 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1783] = heapMem[localMem[1677]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3952;
      end

       3952 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1783]] = 1;
              ip = 3953;
      end

       3953 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1784] = heapMem[localMem[1677]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3954;
      end

       3954 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1784]] = 2;
              ip = 3955;
      end

       3955 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3957;
      end

       3956 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3962;
      end

       3957 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3958;
      end

       3958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1678] = 1;
              updateArrayLength(2, 0, 0);
              ip = 3959;
      end

       3959 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3962;
      end

       3960 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3961;
      end

       3961 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1678] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3962;
      end

       3962 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3963;
      end

       3963 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1678] != 0 ? 3965 : 3964;
      end

       3964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1449] = localMem[1677];
              updateArrayLength(2, 0, 0);
              ip = 3965;
      end

       3965 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3966;
      end

       3966 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3967;
      end

       3967 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1557] = localMem[1557] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3968;
      end

       3968 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3470;
      end

       3969 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3970;
      end

       3970 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
            ip = 3971;
      end

       3971 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3972;
      end

       3972 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3973;
      end

       3973 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3974;
      end

       3974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1785] = heapMem[localMem[1426]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3975;
      end

       3975 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1786] = heapMem[localMem[1426]*6 + 1];
              updateArrayLength(2, 0, 0);
              ip = 3976;
      end

       3976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1787] = heapMem[localMem[1426]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3977;
      end

       3977 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1786] != 1 ? 3981 : 3978;
      end

       3978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1788] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3979;
      end

       3979 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1788]*6 + localMem[1787]] = 44;
              updateArrayLength(1, localMem[1788], localMem[1787]);
              ip = 3980;
      end

       3980 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4227;
      end

       3981 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3982;
      end

       3982 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1786] != 2 ? 3990 : 3983;
      end

       3983 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1789] = localMem[1787] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3984;
      end

       3984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1790] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3985;
      end

       3985 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1790] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1789], localMem[1790], arraySizes[localMem[1790]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1789] && i <= arraySizes[localMem[1790]]) begin
                  heapMem[NArea * localMem[1790] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1790] + localMem[1789]] = 4;                                    // Insert new value
              arraySizes[localMem[1790]] = arraySizes[localMem[1790]] + 1;                              // Increase array size
              ip = 3986;
      end

       3986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1791] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3987;
      end

       3987 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1791] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1789], localMem[1791], arraySizes[localMem[1791]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1789] && i <= arraySizes[localMem[1791]]) begin
                  heapMem[NArea * localMem[1791] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1791] + localMem[1789]] = 44;                                    // Insert new value
              arraySizes[localMem[1791]] = arraySizes[localMem[1791]] + 1;                              // Increase array size
              ip = 3988;
      end

       3988 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1785]*6 + 0] = heapMem[localMem[1785]*6 + 0] + 1;
              updateArrayLength(1, localMem[1785], 0);
              ip = 3989;
      end

       3989 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3996;
      end

       3990 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3991;
      end

       3991 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1792] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3992;
      end

       3992 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1792] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1787], localMem[1792], arraySizes[localMem[1792]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1787] && i <= arraySizes[localMem[1792]]) begin
                  heapMem[NArea * localMem[1792] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1792] + localMem[1787]] = 4;                                    // Insert new value
              arraySizes[localMem[1792]] = arraySizes[localMem[1792]] + 1;                              // Increase array size
              ip = 3993;
      end

       3993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1793] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3994;
      end

       3994 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1793] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1787], localMem[1793], arraySizes[localMem[1793]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1787] && i <= arraySizes[localMem[1793]]) begin
                  heapMem[NArea * localMem[1793] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1793] + localMem[1787]] = 44;                                    // Insert new value
              arraySizes[localMem[1793]] = arraySizes[localMem[1793]] + 1;                              // Increase array size
              ip = 3995;
      end

       3995 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1785]*6 + 0] = heapMem[localMem[1785]*6 + 0] + 1;
              updateArrayLength(1, localMem[1785], 0);
              ip = 3996;
      end

       3996 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3997;
      end

       3997 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 3998;
      end

       3998 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3999;
      end

       3999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1795] = heapMem[localMem[1785]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4000;
      end

       4000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1796] = heapMem[localMem[1785]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4001;
      end

       4001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1797] = heapMem[localMem[1796]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4002;
      end

       4002 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1795] <  localMem[1797] ? 4222 : 4003;
      end

       4003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1798] = localMem[1797];
              updateArrayLength(2, 0, 0);
              ip = 4004;
      end

       4004 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1798] = localMem[1798] >> 1;
              ip = 4005;
      end

       4005 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1799] = localMem[1798] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4006;
      end

       4006 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1800] = heapMem[localMem[1785]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4007;
      end

       4007 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1800] == 0 ? 4104 : 4008;
      end

       4008 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1801] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1801] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1801]] = 0;
              ip = 4009;
      end

       4009 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 0] = localMem[1798];
              updateArrayLength(1, localMem[1801], 0);
              ip = 4010;
      end

       4010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 2] = 0;
              updateArrayLength(1, localMem[1801], 2);
              ip = 4011;
      end

       4011 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1802] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1802] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1802]] = 0;
              ip = 4012;
      end

       4012 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 4] = localMem[1802];
              updateArrayLength(1, localMem[1801], 4);
              ip = 4013;
      end

       4013 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1803] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1803] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1803]] = 0;
              ip = 4014;
      end

       4014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 5] = localMem[1803];
              updateArrayLength(1, localMem[1801], 5);
              ip = 4015;
      end

       4015 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 6] = 0;
              updateArrayLength(1, localMem[1801], 6);
              ip = 4016;
      end

       4016 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 3] = localMem[1796];
              updateArrayLength(1, localMem[1801], 3);
              ip = 4017;
      end

       4017 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1796]*6 + 1] = heapMem[localMem[1796]*6 + 1] + 1;
              updateArrayLength(1, localMem[1796], 1);
              ip = 4018;
      end

       4018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 1] = heapMem[localMem[1796]*6 + 1];
              updateArrayLength(1, localMem[1801], 1);
              ip = 4019;
      end

       4019 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1804] = !heapMem[localMem[1785]*6 + 6];
              ip = 4020;
      end

       4020 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1804] != 0 ? 4049 : 4021;
      end

       4021 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1805] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1805] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1805]] = 0;
              ip = 4022;
      end

       4022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 6] = localMem[1805];
              updateArrayLength(1, localMem[1801], 6);
              ip = 4023;
      end

       4023 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1806] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4024;
      end

       4024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1807] = heapMem[localMem[1801]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4025;
      end

       4025 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1807] + 0 + i] = heapMem[NArea * localMem[1806] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1807], 0 + i);
                end
              end
              ip = 4026;
      end

       4026 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1808] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4027;
      end

       4027 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1809] = heapMem[localMem[1801]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4028;
      end

       4028 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1809] + 0 + i] = heapMem[NArea * localMem[1808] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1809], 0 + i);
                end
              end
              ip = 4029;
      end

       4029 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1810] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4030;
      end

       4030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1811] = heapMem[localMem[1801]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4031;
      end

       4031 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1812] = localMem[1798] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4032;
      end

       4032 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1812]) begin
                  heapMem[NArea * localMem[1811] + 0 + i] = heapMem[NArea * localMem[1810] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1811], 0 + i);
                end
              end
              ip = 4033;
      end

       4033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1813] = heapMem[localMem[1801]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4034;
      end

       4034 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1814] = localMem[1813] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4035;
      end

       4035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1815] = heapMem[localMem[1801]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4036;
      end

       4036 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4037;
      end

       4037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1816] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4038;
      end

       4038 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4039;
      end

       4039 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1816] >= localMem[1814] ? 4045 : 4040;
      end

       4040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1817] = heapMem[localMem[1815]*6 + localMem[1816]];
              updateArrayLength(2, 0, 0);
              ip = 4041;
      end

       4041 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1817]*6 + 2] = localMem[1801];
              updateArrayLength(1, localMem[1817], 2);
              ip = 4042;
      end

       4042 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4043;
      end

       4043 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1816] = localMem[1816] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4044;
      end

       4044 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4038;
      end

       4045 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4046;
      end

       4046 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1818] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4047;
      end

       4047 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1818]] = localMem[1799];
              ip = 4048;
      end

       4048 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4056;
      end

       4049 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4050;
      end

       4050 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1819] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4051;
      end

       4051 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1820] = heapMem[localMem[1801]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4052;
      end

       4052 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1820] + 0 + i] = heapMem[NArea * localMem[1819] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1820], 0 + i);
                end
              end
              ip = 4053;
      end

       4053 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1821] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4054;
      end

       4054 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1822] = heapMem[localMem[1801]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4055;
      end

       4055 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1822] + 0 + i] = heapMem[NArea * localMem[1821] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1822], 0 + i);
                end
              end
              ip = 4056;
      end

       4056 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4057;
      end

       4057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1785]*6 + 0] = localMem[1798];
              updateArrayLength(1, localMem[1785], 0);
              ip = 4058;
      end

       4058 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1801]*6 + 2] = localMem[1800];
              updateArrayLength(1, localMem[1801], 2);
              ip = 4059;
      end

       4059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1823] = heapMem[localMem[1800]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4060;
      end

       4060 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1824] = heapMem[localMem[1800]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4061;
      end

       4061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1825] = heapMem[localMem[1824]*6 + localMem[1823]];
              updateArrayLength(2, 0, 0);
              ip = 4062;
      end

       4062 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1825] != localMem[1785] ? 4081 : 4063;
      end

       4063 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1826] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4064;
      end

       4064 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1827] = heapMem[localMem[1826]*6 + localMem[1798]];
              updateArrayLength(2, 0, 0);
              ip = 4065;
      end

       4065 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1828] = heapMem[localMem[1800]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4066;
      end

       4066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1828]*6 + localMem[1823]] = localMem[1827];
              updateArrayLength(1, localMem[1828], localMem[1823]);
              ip = 4067;
      end

       4067 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1829] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4068;
      end

       4068 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1830] = heapMem[localMem[1829]*6 + localMem[1798]];
              updateArrayLength(2, 0, 0);
              ip = 4069;
      end

       4069 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1831] = heapMem[localMem[1800]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4070;
      end

       4070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1831]*6 + localMem[1823]] = localMem[1830];
              updateArrayLength(1, localMem[1831], localMem[1823]);
              ip = 4071;
      end

       4071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1832] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4072;
      end

       4072 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1832]] = localMem[1798];
              ip = 4073;
      end

       4073 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1833] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4074;
      end

       4074 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1833]] = localMem[1798];
              ip = 4075;
      end

       4075 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1834] = localMem[1823] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4076;
      end

       4076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1800]*6 + 0] = localMem[1834];
              updateArrayLength(1, localMem[1800], 0);
              ip = 4077;
      end

       4077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1835] = heapMem[localMem[1800]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4078;
      end

       4078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1835]*6 + localMem[1834]] = localMem[1801];
              updateArrayLength(1, localMem[1835], localMem[1834]);
              ip = 4079;
      end

       4079 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4219;
      end

       4080 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4103;
      end

       4081 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4082;
      end

       4082 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 4083;
      end

       4083 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1836] = heapMem[localMem[1800]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4084;
      end

       4084 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1837] = 0; k = arraySizes[localMem[1836]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1836] * NArea + i] == localMem[1785]) localMem[1837] = i + 1;
              end
              ip = 4085;
      end

       4085 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1837] = localMem[1837] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4086;
      end

       4086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1838] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4087;
      end

       4087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1839] = heapMem[localMem[1838]*6 + localMem[1798]];
              updateArrayLength(2, 0, 0);
              ip = 4088;
      end

       4088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1840] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4089;
      end

       4089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1841] = heapMem[localMem[1840]*6 + localMem[1798]];
              updateArrayLength(2, 0, 0);
              ip = 4090;
      end

       4090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1842] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4091;
      end

       4091 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1842]] = localMem[1798];
              ip = 4092;
      end

       4092 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1843] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4093;
      end

       4093 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1843]] = localMem[1798];
              ip = 4094;
      end

       4094 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1844] = heapMem[localMem[1800]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4095;
      end

       4095 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1844] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1837], localMem[1844], arraySizes[localMem[1844]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1837] && i <= arraySizes[localMem[1844]]) begin
                  heapMem[NArea * localMem[1844] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1844] + localMem[1837]] = localMem[1839];                                    // Insert new value
              arraySizes[localMem[1844]] = arraySizes[localMem[1844]] + 1;                              // Increase array size
              ip = 4096;
      end

       4096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1845] = heapMem[localMem[1800]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4097;
      end

       4097 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1845] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1837], localMem[1845], arraySizes[localMem[1845]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1837] && i <= arraySizes[localMem[1845]]) begin
                  heapMem[NArea * localMem[1845] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1845] + localMem[1837]] = localMem[1841];                                    // Insert new value
              arraySizes[localMem[1845]] = arraySizes[localMem[1845]] + 1;                              // Increase array size
              ip = 4098;
      end

       4098 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1846] = heapMem[localMem[1800]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4099;
      end

       4099 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1847] = localMem[1837] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4100;
      end

       4100 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1846] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1847], localMem[1846], arraySizes[localMem[1846]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1847] && i <= arraySizes[localMem[1846]]) begin
                  heapMem[NArea * localMem[1846] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1846] + localMem[1847]] = localMem[1801];                                    // Insert new value
              arraySizes[localMem[1846]] = arraySizes[localMem[1846]] + 1;                              // Increase array size
              ip = 4101;
      end

       4101 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1800]*6 + 0] = heapMem[localMem[1800]*6 + 0] + 1;
              updateArrayLength(1, localMem[1800], 0);
              ip = 4102;
      end

       4102 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4219;
      end

       4103 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4104;
      end

       4104 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4105;
      end

       4105 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1848] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1848] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1848]] = 0;
              ip = 4106;
      end

       4106 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 0] = localMem[1798];
              updateArrayLength(1, localMem[1848], 0);
              ip = 4107;
      end

       4107 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 2] = 0;
              updateArrayLength(1, localMem[1848], 2);
              ip = 4108;
      end

       4108 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1849] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1849] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1849]] = 0;
              ip = 4109;
      end

       4109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 4] = localMem[1849];
              updateArrayLength(1, localMem[1848], 4);
              ip = 4110;
      end

       4110 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1850] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1850] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1850]] = 0;
              ip = 4111;
      end

       4111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 5] = localMem[1850];
              updateArrayLength(1, localMem[1848], 5);
              ip = 4112;
      end

       4112 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 6] = 0;
              updateArrayLength(1, localMem[1848], 6);
              ip = 4113;
      end

       4113 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 3] = localMem[1796];
              updateArrayLength(1, localMem[1848], 3);
              ip = 4114;
      end

       4114 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1796]*6 + 1] = heapMem[localMem[1796]*6 + 1] + 1;
              updateArrayLength(1, localMem[1796], 1);
              ip = 4115;
      end

       4115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 1] = heapMem[localMem[1796]*6 + 1];
              updateArrayLength(1, localMem[1848], 1);
              ip = 4116;
      end

       4116 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1851] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1851] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1851]] = 0;
              ip = 4117;
      end

       4117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 0] = localMem[1798];
              updateArrayLength(1, localMem[1851], 0);
              ip = 4118;
      end

       4118 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 2] = 0;
              updateArrayLength(1, localMem[1851], 2);
              ip = 4119;
      end

       4119 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1852] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1852] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1852]] = 0;
              ip = 4120;
      end

       4120 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 4] = localMem[1852];
              updateArrayLength(1, localMem[1851], 4);
              ip = 4121;
      end

       4121 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1853] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1853] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1853]] = 0;
              ip = 4122;
      end

       4122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 5] = localMem[1853];
              updateArrayLength(1, localMem[1851], 5);
              ip = 4123;
      end

       4123 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 6] = 0;
              updateArrayLength(1, localMem[1851], 6);
              ip = 4124;
      end

       4124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 3] = localMem[1796];
              updateArrayLength(1, localMem[1851], 3);
              ip = 4125;
      end

       4125 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1796]*6 + 1] = heapMem[localMem[1796]*6 + 1] + 1;
              updateArrayLength(1, localMem[1796], 1);
              ip = 4126;
      end

       4126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 1] = heapMem[localMem[1796]*6 + 1];
              updateArrayLength(1, localMem[1851], 1);
              ip = 4127;
      end

       4127 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1854] = !heapMem[localMem[1785]*6 + 6];
              ip = 4128;
      end

       4128 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1854] != 0 ? 4180 : 4129;
      end

       4129 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1855] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1855] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1855]] = 0;
              ip = 4130;
      end

       4130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 6] = localMem[1855];
              updateArrayLength(1, localMem[1848], 6);
              ip = 4131;
      end

       4131 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1856] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1856] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1856]] = 0;
              ip = 4132;
      end

       4132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 6] = localMem[1856];
              updateArrayLength(1, localMem[1851], 6);
              ip = 4133;
      end

       4133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1857] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4134;
      end

       4134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1858] = heapMem[localMem[1848]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4135;
      end

       4135 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1858] + 0 + i] = heapMem[NArea * localMem[1857] + 0 + i];
                  updateArrayLength(1, localMem[1858], 0 + i);
                end
              end
              ip = 4136;
      end

       4136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1859] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4137;
      end

       4137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1860] = heapMem[localMem[1848]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4138;
      end

       4138 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1860] + 0 + i] = heapMem[NArea * localMem[1859] + 0 + i];
                  updateArrayLength(1, localMem[1860], 0 + i);
                end
              end
              ip = 4139;
      end

       4139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1861] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4140;
      end

       4140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1862] = heapMem[localMem[1848]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4141;
      end

       4141 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1863] = localMem[1798] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4142;
      end

       4142 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1863]) begin
                  heapMem[NArea * localMem[1862] + 0 + i] = heapMem[NArea * localMem[1861] + 0 + i];
                  updateArrayLength(1, localMem[1862], 0 + i);
                end
              end
              ip = 4143;
      end

       4143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1864] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4144;
      end

       4144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1865] = heapMem[localMem[1851]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4145;
      end

       4145 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1865] + 0 + i] = heapMem[NArea * localMem[1864] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1865], 0 + i);
                end
              end
              ip = 4146;
      end

       4146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1866] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4147;
      end

       4147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1867] = heapMem[localMem[1851]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4148;
      end

       4148 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1867] + 0 + i] = heapMem[NArea * localMem[1866] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1867], 0 + i);
                end
              end
              ip = 4149;
      end

       4149 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1868] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4150;
      end

       4150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1869] = heapMem[localMem[1851]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4151;
      end

       4151 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1870] = localMem[1798] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4152;
      end

       4152 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1870]) begin
                  heapMem[NArea * localMem[1869] + 0 + i] = heapMem[NArea * localMem[1868] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1869], 0 + i);
                end
              end
              ip = 4153;
      end

       4153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1871] = heapMem[localMem[1848]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4154;
      end

       4154 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1872] = localMem[1871] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4155;
      end

       4155 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1873] = heapMem[localMem[1848]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4156;
      end

       4156 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4157;
      end

       4157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1874] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4158;
      end

       4158 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4159;
      end

       4159 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1874] >= localMem[1872] ? 4165 : 4160;
      end

       4160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1875] = heapMem[localMem[1873]*6 + localMem[1874]];
              updateArrayLength(2, 0, 0);
              ip = 4161;
      end

       4161 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1875]*6 + 2] = localMem[1848];
              updateArrayLength(1, localMem[1875], 2);
              ip = 4162;
      end

       4162 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4163;
      end

       4163 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1874] = localMem[1874] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4164;
      end

       4164 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4158;
      end

       4165 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4166;
      end

       4166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1876] = heapMem[localMem[1851]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4167;
      end

       4167 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1877] = localMem[1876] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4168;
      end

       4168 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1878] = heapMem[localMem[1851]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4169;
      end

       4169 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4170;
      end

       4170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1879] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4171;
      end

       4171 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4172;
      end

       4172 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1879] >= localMem[1877] ? 4178 : 4173;
      end

       4173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1880] = heapMem[localMem[1878]*6 + localMem[1879]];
              updateArrayLength(2, 0, 0);
              ip = 4174;
      end

       4174 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1880]*6 + 2] = localMem[1851];
              updateArrayLength(1, localMem[1880], 2);
              ip = 4175;
      end

       4175 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4176;
      end

       4176 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1879] = localMem[1879] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4177;
      end

       4177 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4171;
      end

       4178 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4179;
      end

       4179 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4195;
      end

       4180 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4181;
      end

       4181 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1881] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1881] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1881]] = 0;
              ip = 4182;
      end

       4182 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1785]*6 + 6] = localMem[1881];
              updateArrayLength(1, localMem[1785], 6);
              ip = 4183;
      end

       4183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1882] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4184;
      end

       4184 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1883] = heapMem[localMem[1848]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4185;
      end

       4185 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1883] + 0 + i] = heapMem[NArea * localMem[1882] + 0 + i];
                  updateArrayLength(1, localMem[1883], 0 + i);
                end
              end
              ip = 4186;
      end

       4186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1884] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4187;
      end

       4187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1885] = heapMem[localMem[1848]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4188;
      end

       4188 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1885] + 0 + i] = heapMem[NArea * localMem[1884] + 0 + i];
                  updateArrayLength(1, localMem[1885], 0 + i);
                end
              end
              ip = 4189;
      end

       4189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1886] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4190;
      end

       4190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1887] = heapMem[localMem[1851]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4191;
      end

       4191 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1887] + 0 + i] = heapMem[NArea * localMem[1886] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1887], 0 + i);
                end
              end
              ip = 4192;
      end

       4192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1888] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4193;
      end

       4193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1889] = heapMem[localMem[1851]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4194;
      end

       4194 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1798]) begin
                  heapMem[NArea * localMem[1889] + 0 + i] = heapMem[NArea * localMem[1888] + localMem[1799] + i];
                  updateArrayLength(1, localMem[1889], 0 + i);
                end
              end
              ip = 4195;
      end

       4195 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4196;
      end

       4196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1848]*6 + 2] = localMem[1785];
              updateArrayLength(1, localMem[1848], 2);
              ip = 4197;
      end

       4197 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1851]*6 + 2] = localMem[1785];
              updateArrayLength(1, localMem[1851], 2);
              ip = 4198;
      end

       4198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1890] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4199;
      end

       4199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1891] = heapMem[localMem[1890]*6 + localMem[1798]];
              updateArrayLength(2, 0, 0);
              ip = 4200;
      end

       4200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1892] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4201;
      end

       4201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1893] = heapMem[localMem[1892]*6 + localMem[1798]];
              updateArrayLength(2, 0, 0);
              ip = 4202;
      end

       4202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1894] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4203;
      end

       4203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1894]*6 + 0] = localMem[1891];
              updateArrayLength(1, localMem[1894], 0);
              ip = 4204;
      end

       4204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1895] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4205;
      end

       4205 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1895]*6 + 0] = localMem[1893];
              updateArrayLength(1, localMem[1895], 0);
              ip = 4206;
      end

       4206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1896] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4207;
      end

       4207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1896]*6 + 0] = localMem[1848];
              updateArrayLength(1, localMem[1896], 0);
              ip = 4208;
      end

       4208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1897] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4209;
      end

       4209 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1897]*6 + 1] = localMem[1851];
              updateArrayLength(1, localMem[1897], 1);
              ip = 4210;
      end

       4210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1785]*6 + 0] = 1;
              updateArrayLength(1, localMem[1785], 0);
              ip = 4211;
      end

       4211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1898] = heapMem[localMem[1785]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4212;
      end

       4212 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1898]] = 1;
              ip = 4213;
      end

       4213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1899] = heapMem[localMem[1785]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4214;
      end

       4214 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1899]] = 1;
              ip = 4215;
      end

       4215 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1900] = heapMem[localMem[1785]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4216;
      end

       4216 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1900]] = 2;
              ip = 4217;
      end

       4217 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4219;
      end

       4218 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4224;
      end

       4219 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4220;
      end

       4220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1794] = 1;
              updateArrayLength(2, 0, 0);
              ip = 4221;
      end

       4221 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4224;
      end

       4222 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4223;
      end

       4223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1794] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4224;
      end

       4224 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4225;
      end

       4225 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4226;
      end

       4226 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4227;
      end

       4227 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4228;
      end

       4228 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[1426]] = 0;
              freedArrays[freedArraysTop] = localMem[1426];
              freedArraysTop = freedArraysTop + 1;
              ip = 4229;
      end

       4229 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1901] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1901] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1901]] = 0;
              ip = 4230;
      end

       4230 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4231;
      end

       4231 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1902] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4232;
      end

       4232 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1902] != 0 ? 4255 : 4233;
      end

       4233 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1903] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1903] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1903]] = 0;
              ip = 4234;
      end

       4234 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 0] = 1;
              updateArrayLength(1, localMem[1903], 0);
              ip = 4235;
      end

       4235 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 2] = 0;
              updateArrayLength(1, localMem[1903], 2);
              ip = 4236;
      end

       4236 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1904] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1904] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1904]] = 0;
              ip = 4237;
      end

       4237 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 4] = localMem[1904];
              updateArrayLength(1, localMem[1903], 4);
              ip = 4238;
      end

       4238 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1905] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1905] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1905]] = 0;
              ip = 4239;
      end

       4239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 5] = localMem[1905];
              updateArrayLength(1, localMem[1903], 5);
              ip = 4240;
      end

       4240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 6] = 0;
              updateArrayLength(1, localMem[1903], 6);
              ip = 4241;
      end

       4241 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 3] = localMem[0];
              updateArrayLength(1, localMem[1903], 3);
              ip = 4242;
      end

       4242 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = heapMem[localMem[0]*6 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 4243;
      end

       4243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1903]*6 + 1] = heapMem[localMem[0]*6 + 1];
              updateArrayLength(1, localMem[1903], 1);
              ip = 4244;
      end

       4244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1906] = heapMem[localMem[1903]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4245;
      end

       4245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1906]*6 + 0] = 5;
              updateArrayLength(1, localMem[1906], 0);
              ip = 4246;
      end

       4246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1907] = heapMem[localMem[1903]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4247;
      end

       4247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1907]*6 + 0] = 55;
              updateArrayLength(1, localMem[1907], 0);
              ip = 4248;
      end

       4248 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 4249;
      end

       4249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = localMem[1903];
              updateArrayLength(1, localMem[0], 3);
              ip = 4250;
      end

       4250 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1908] = heapMem[localMem[1903]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4251;
      end

       4251 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1908]] = 1;
              ip = 4252;
      end

       4252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1909] = heapMem[localMem[1903]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4253;
      end

       4253 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1909]] = 1;
              ip = 4254;
      end

       4254 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5283;
      end

       4255 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4256;
      end

       4256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1910] = heapMem[localMem[1902]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4257;
      end

       4257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1911] = heapMem[localMem[0]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4258;
      end

       4258 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1910] >= localMem[1911] ? 4294 : 4259;
      end

       4259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1912] = heapMem[localMem[1902]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4260;
      end

       4260 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1912] != 0 ? 4293 : 4261;
      end

       4261 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1913] = !heapMem[localMem[1902]*6 + 6];
              ip = 4262;
      end

       4262 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1913] == 0 ? 4292 : 4263;
      end

       4263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1914] = heapMem[localMem[1902]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4264;
      end

       4264 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1915] = 0; k = arraySizes[localMem[1914]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1914] * NArea + i] == 5) localMem[1915] = i + 1;
              end
              ip = 4265;
      end

       4265 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1915] == 0 ? 4270 : 4266;
      end

       4266 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1915] = localMem[1915] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4267;
      end

       4267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1916] = heapMem[localMem[1902]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4268;
      end

       4268 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1916]*6 + localMem[1915]] = 55;
              updateArrayLength(1, localMem[1916], localMem[1915]);
              ip = 4269;
      end

       4269 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5283;
      end

       4270 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4271;
      end

       4271 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1914]] = localMem[1910];
              ip = 4272;
      end

       4272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1917] = heapMem[localMem[1902]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4273;
      end

       4273 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1917]] = localMem[1910];
              ip = 4274;
      end

       4274 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[1914]];
//$display("AAAAA k=%d  source2=%d", k, 5);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[1914] * NArea + i]);
                if (i < k && heapMem[localMem[1914] * NArea + i] > 5) j = j + 1;
              end
              localMem[1918] = j;
              ip = 4275;
      end

       4275 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1918] != 0 ? 4283 : 4276;
      end

       4276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1919] = heapMem[localMem[1902]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4277;
      end

       4277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1919]*6 + localMem[1910]] = 5;
              updateArrayLength(1, localMem[1919], localMem[1910]);
              ip = 4278;
      end

       4278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1920] = heapMem[localMem[1902]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4279;
      end

       4279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1920]*6 + localMem[1910]] = 55;
              updateArrayLength(1, localMem[1920], localMem[1910]);
              ip = 4280;
      end

       4280 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1902]*6 + 0] = localMem[1910] + 1;
              updateArrayLength(1, localMem[1902], 0);
              ip = 4281;
      end

       4281 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 4282;
      end

       4282 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5283;
      end

       4283 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4284;
      end

       4284 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[1914]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1914] * NArea + i] < 5) j = j + 1;
              end
              localMem[1921] = j;
              ip = 4285;
      end

       4285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1922] = heapMem[localMem[1902]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4286;
      end

       4286 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1922] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1921], localMem[1922], arraySizes[localMem[1922]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1921] && i <= arraySizes[localMem[1922]]) begin
                  heapMem[NArea * localMem[1922] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1922] + localMem[1921]] = 5;                                    // Insert new value
              arraySizes[localMem[1922]] = arraySizes[localMem[1922]] + 1;                              // Increase array size
              ip = 4287;
      end

       4287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1923] = heapMem[localMem[1902]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4288;
      end

       4288 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1923] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1921], localMem[1923], arraySizes[localMem[1923]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1921] && i <= arraySizes[localMem[1923]]) begin
                  heapMem[NArea * localMem[1923] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1923] + localMem[1921]] = 55;                                    // Insert new value
              arraySizes[localMem[1923]] = arraySizes[localMem[1923]] + 1;                              // Increase array size
              ip = 4289;
      end

       4289 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1902]*6 + 0] = heapMem[localMem[1902]*6 + 0] + 1;
              updateArrayLength(1, localMem[1902], 0);
              ip = 4290;
      end

       4290 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 4291;
      end

       4291 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5283;
      end

       4292 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4293;
      end

       4293 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4294;
      end

       4294 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4295;
      end

       4295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1924] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4296;
      end

       4296 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4297;
      end

       4297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1926] = heapMem[localMem[1924]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4298;
      end

       4298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1927] = heapMem[localMem[1924]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4299;
      end

       4299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1928] = heapMem[localMem[1927]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4300;
      end

       4300 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1926] <  localMem[1928] ? 4520 : 4301;
      end

       4301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1929] = localMem[1928];
              updateArrayLength(2, 0, 0);
              ip = 4302;
      end

       4302 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1929] = localMem[1929] >> 1;
              ip = 4303;
      end

       4303 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1930] = localMem[1929] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4304;
      end

       4304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1931] = heapMem[localMem[1924]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4305;
      end

       4305 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1931] == 0 ? 4402 : 4306;
      end

       4306 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1932] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1932] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1932]] = 0;
              ip = 4307;
      end

       4307 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 0] = localMem[1929];
              updateArrayLength(1, localMem[1932], 0);
              ip = 4308;
      end

       4308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 2] = 0;
              updateArrayLength(1, localMem[1932], 2);
              ip = 4309;
      end

       4309 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1933] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1933] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1933]] = 0;
              ip = 4310;
      end

       4310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 4] = localMem[1933];
              updateArrayLength(1, localMem[1932], 4);
              ip = 4311;
      end

       4311 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1934] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1934] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1934]] = 0;
              ip = 4312;
      end

       4312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 5] = localMem[1934];
              updateArrayLength(1, localMem[1932], 5);
              ip = 4313;
      end

       4313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 6] = 0;
              updateArrayLength(1, localMem[1932], 6);
              ip = 4314;
      end

       4314 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 3] = localMem[1927];
              updateArrayLength(1, localMem[1932], 3);
              ip = 4315;
      end

       4315 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1927]*6 + 1] = heapMem[localMem[1927]*6 + 1] + 1;
              updateArrayLength(1, localMem[1927], 1);
              ip = 4316;
      end

       4316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 1] = heapMem[localMem[1927]*6 + 1];
              updateArrayLength(1, localMem[1932], 1);
              ip = 4317;
      end

       4317 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1935] = !heapMem[localMem[1924]*6 + 6];
              ip = 4318;
      end

       4318 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1935] != 0 ? 4347 : 4319;
      end

       4319 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1936] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1936] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1936]] = 0;
              ip = 4320;
      end

       4320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 6] = localMem[1936];
              updateArrayLength(1, localMem[1932], 6);
              ip = 4321;
      end

       4321 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1937] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4322;
      end

       4322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1938] = heapMem[localMem[1932]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4323;
      end

       4323 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1938] + 0 + i] = heapMem[NArea * localMem[1937] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1938], 0 + i);
                end
              end
              ip = 4324;
      end

       4324 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1939] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4325;
      end

       4325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1940] = heapMem[localMem[1932]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4326;
      end

       4326 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1940] + 0 + i] = heapMem[NArea * localMem[1939] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1940], 0 + i);
                end
              end
              ip = 4327;
      end

       4327 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1941] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4328;
      end

       4328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1942] = heapMem[localMem[1932]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4329;
      end

       4329 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1943] = localMem[1929] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4330;
      end

       4330 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1943]) begin
                  heapMem[NArea * localMem[1942] + 0 + i] = heapMem[NArea * localMem[1941] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1942], 0 + i);
                end
              end
              ip = 4331;
      end

       4331 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1944] = heapMem[localMem[1932]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4332;
      end

       4332 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1945] = localMem[1944] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4333;
      end

       4333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1946] = heapMem[localMem[1932]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4334;
      end

       4334 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4335;
      end

       4335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1947] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4336;
      end

       4336 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4337;
      end

       4337 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1947] >= localMem[1945] ? 4343 : 4338;
      end

       4338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1948] = heapMem[localMem[1946]*6 + localMem[1947]];
              updateArrayLength(2, 0, 0);
              ip = 4339;
      end

       4339 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1948]*6 + 2] = localMem[1932];
              updateArrayLength(1, localMem[1948], 2);
              ip = 4340;
      end

       4340 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4341;
      end

       4341 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1947] = localMem[1947] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4342;
      end

       4342 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4336;
      end

       4343 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4344;
      end

       4344 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1949] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4345;
      end

       4345 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1949]] = localMem[1930];
              ip = 4346;
      end

       4346 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4354;
      end

       4347 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4348;
      end

       4348 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1950] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4349;
      end

       4349 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1951] = heapMem[localMem[1932]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4350;
      end

       4350 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1951] + 0 + i] = heapMem[NArea * localMem[1950] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1951], 0 + i);
                end
              end
              ip = 4351;
      end

       4351 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1952] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4352;
      end

       4352 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1953] = heapMem[localMem[1932]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4353;
      end

       4353 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1953] + 0 + i] = heapMem[NArea * localMem[1952] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1953], 0 + i);
                end
              end
              ip = 4354;
      end

       4354 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4355;
      end

       4355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1924]*6 + 0] = localMem[1929];
              updateArrayLength(1, localMem[1924], 0);
              ip = 4356;
      end

       4356 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1932]*6 + 2] = localMem[1931];
              updateArrayLength(1, localMem[1932], 2);
              ip = 4357;
      end

       4357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1954] = heapMem[localMem[1931]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4358;
      end

       4358 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1955] = heapMem[localMem[1931]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4359;
      end

       4359 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1956] = heapMem[localMem[1955]*6 + localMem[1954]];
              updateArrayLength(2, 0, 0);
              ip = 4360;
      end

       4360 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1956] != localMem[1924] ? 4379 : 4361;
      end

       4361 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1957] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4362;
      end

       4362 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1958] = heapMem[localMem[1957]*6 + localMem[1929]];
              updateArrayLength(2, 0, 0);
              ip = 4363;
      end

       4363 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1959] = heapMem[localMem[1931]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4364;
      end

       4364 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1959]*6 + localMem[1954]] = localMem[1958];
              updateArrayLength(1, localMem[1959], localMem[1954]);
              ip = 4365;
      end

       4365 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1960] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4366;
      end

       4366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1961] = heapMem[localMem[1960]*6 + localMem[1929]];
              updateArrayLength(2, 0, 0);
              ip = 4367;
      end

       4367 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1962] = heapMem[localMem[1931]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4368;
      end

       4368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1962]*6 + localMem[1954]] = localMem[1961];
              updateArrayLength(1, localMem[1962], localMem[1954]);
              ip = 4369;
      end

       4369 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1963] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4370;
      end

       4370 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1963]] = localMem[1929];
              ip = 4371;
      end

       4371 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1964] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4372;
      end

       4372 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1964]] = localMem[1929];
              ip = 4373;
      end

       4373 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1965] = localMem[1954] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4374;
      end

       4374 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1931]*6 + 0] = localMem[1965];
              updateArrayLength(1, localMem[1931], 0);
              ip = 4375;
      end

       4375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1966] = heapMem[localMem[1931]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4376;
      end

       4376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1966]*6 + localMem[1965]] = localMem[1932];
              updateArrayLength(1, localMem[1966], localMem[1965]);
              ip = 4377;
      end

       4377 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4517;
      end

       4378 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4401;
      end

       4379 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4380;
      end

       4380 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 4381;
      end

       4381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1967] = heapMem[localMem[1931]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4382;
      end

       4382 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[1968] = 0; k = arraySizes[localMem[1967]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[1967] * NArea + i] == localMem[1924]) localMem[1968] = i + 1;
              end
              ip = 4383;
      end

       4383 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1968] = localMem[1968] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4384;
      end

       4384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1969] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4385;
      end

       4385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1970] = heapMem[localMem[1969]*6 + localMem[1929]];
              updateArrayLength(2, 0, 0);
              ip = 4386;
      end

       4386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1971] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4387;
      end

       4387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1972] = heapMem[localMem[1971]*6 + localMem[1929]];
              updateArrayLength(2, 0, 0);
              ip = 4388;
      end

       4388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1973] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4389;
      end

       4389 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1973]] = localMem[1929];
              ip = 4390;
      end

       4390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1974] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4391;
      end

       4391 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1974]] = localMem[1929];
              ip = 4392;
      end

       4392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1975] = heapMem[localMem[1931]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4393;
      end

       4393 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1975] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1968], localMem[1975], arraySizes[localMem[1975]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1968] && i <= arraySizes[localMem[1975]]) begin
                  heapMem[NArea * localMem[1975] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1975] + localMem[1968]] = localMem[1970];                                    // Insert new value
              arraySizes[localMem[1975]] = arraySizes[localMem[1975]] + 1;                              // Increase array size
              ip = 4394;
      end

       4394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1976] = heapMem[localMem[1931]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4395;
      end

       4395 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1976] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1968], localMem[1976], arraySizes[localMem[1976]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1968] && i <= arraySizes[localMem[1976]]) begin
                  heapMem[NArea * localMem[1976] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1976] + localMem[1968]] = localMem[1972];                                    // Insert new value
              arraySizes[localMem[1976]] = arraySizes[localMem[1976]] + 1;                              // Increase array size
              ip = 4396;
      end

       4396 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1977] = heapMem[localMem[1931]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4397;
      end

       4397 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1978] = localMem[1968] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4398;
      end

       4398 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1977] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1978], localMem[1977], arraySizes[localMem[1977]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1978] && i <= arraySizes[localMem[1977]]) begin
                  heapMem[NArea * localMem[1977] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1977] + localMem[1978]] = localMem[1932];                                    // Insert new value
              arraySizes[localMem[1977]] = arraySizes[localMem[1977]] + 1;                              // Increase array size
              ip = 4399;
      end

       4399 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1931]*6 + 0] = heapMem[localMem[1931]*6 + 0] + 1;
              updateArrayLength(1, localMem[1931], 0);
              ip = 4400;
      end

       4400 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4517;
      end

       4401 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4402;
      end

       4402 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4403;
      end

       4403 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1979] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1979] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1979]] = 0;
              ip = 4404;
      end

       4404 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 0] = localMem[1929];
              updateArrayLength(1, localMem[1979], 0);
              ip = 4405;
      end

       4405 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 2] = 0;
              updateArrayLength(1, localMem[1979], 2);
              ip = 4406;
      end

       4406 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1980] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1980] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1980]] = 0;
              ip = 4407;
      end

       4407 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 4] = localMem[1980];
              updateArrayLength(1, localMem[1979], 4);
              ip = 4408;
      end

       4408 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1981] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1981] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1981]] = 0;
              ip = 4409;
      end

       4409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 5] = localMem[1981];
              updateArrayLength(1, localMem[1979], 5);
              ip = 4410;
      end

       4410 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 6] = 0;
              updateArrayLength(1, localMem[1979], 6);
              ip = 4411;
      end

       4411 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 3] = localMem[1927];
              updateArrayLength(1, localMem[1979], 3);
              ip = 4412;
      end

       4412 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1927]*6 + 1] = heapMem[localMem[1927]*6 + 1] + 1;
              updateArrayLength(1, localMem[1927], 1);
              ip = 4413;
      end

       4413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 1] = heapMem[localMem[1927]*6 + 1];
              updateArrayLength(1, localMem[1979], 1);
              ip = 4414;
      end

       4414 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1982] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1982] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1982]] = 0;
              ip = 4415;
      end

       4415 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 0] = localMem[1929];
              updateArrayLength(1, localMem[1982], 0);
              ip = 4416;
      end

       4416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 2] = 0;
              updateArrayLength(1, localMem[1982], 2);
              ip = 4417;
      end

       4417 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1983] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1983] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1983]] = 0;
              ip = 4418;
      end

       4418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 4] = localMem[1983];
              updateArrayLength(1, localMem[1982], 4);
              ip = 4419;
      end

       4419 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1984] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1984] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1984]] = 0;
              ip = 4420;
      end

       4420 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 5] = localMem[1984];
              updateArrayLength(1, localMem[1982], 5);
              ip = 4421;
      end

       4421 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 6] = 0;
              updateArrayLength(1, localMem[1982], 6);
              ip = 4422;
      end

       4422 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 3] = localMem[1927];
              updateArrayLength(1, localMem[1982], 3);
              ip = 4423;
      end

       4423 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1927]*6 + 1] = heapMem[localMem[1927]*6 + 1] + 1;
              updateArrayLength(1, localMem[1927], 1);
              ip = 4424;
      end

       4424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 1] = heapMem[localMem[1927]*6 + 1];
              updateArrayLength(1, localMem[1982], 1);
              ip = 4425;
      end

       4425 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1985] = !heapMem[localMem[1924]*6 + 6];
              ip = 4426;
      end

       4426 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1985] != 0 ? 4478 : 4427;
      end

       4427 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1986] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1986] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1986]] = 0;
              ip = 4428;
      end

       4428 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 6] = localMem[1986];
              updateArrayLength(1, localMem[1979], 6);
              ip = 4429;
      end

       4429 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1987] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1987] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1987]] = 0;
              ip = 4430;
      end

       4430 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 6] = localMem[1987];
              updateArrayLength(1, localMem[1982], 6);
              ip = 4431;
      end

       4431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1988] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4432;
      end

       4432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1989] = heapMem[localMem[1979]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4433;
      end

       4433 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1989] + 0 + i] = heapMem[NArea * localMem[1988] + 0 + i];
                  updateArrayLength(1, localMem[1989], 0 + i);
                end
              end
              ip = 4434;
      end

       4434 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1990] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4435;
      end

       4435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1991] = heapMem[localMem[1979]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4436;
      end

       4436 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1991] + 0 + i] = heapMem[NArea * localMem[1990] + 0 + i];
                  updateArrayLength(1, localMem[1991], 0 + i);
                end
              end
              ip = 4437;
      end

       4437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1992] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4438;
      end

       4438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1993] = heapMem[localMem[1979]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4439;
      end

       4439 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1994] = localMem[1929] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4440;
      end

       4440 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1994]) begin
                  heapMem[NArea * localMem[1993] + 0 + i] = heapMem[NArea * localMem[1992] + 0 + i];
                  updateArrayLength(1, localMem[1993], 0 + i);
                end
              end
              ip = 4441;
      end

       4441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1995] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4442;
      end

       4442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1996] = heapMem[localMem[1982]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4443;
      end

       4443 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1996] + 0 + i] = heapMem[NArea * localMem[1995] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1996], 0 + i);
                end
              end
              ip = 4444;
      end

       4444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1997] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4445;
      end

       4445 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1998] = heapMem[localMem[1982]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4446;
      end

       4446 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[1998] + 0 + i] = heapMem[NArea * localMem[1997] + localMem[1930] + i];
                  updateArrayLength(1, localMem[1998], 0 + i);
                end
              end
              ip = 4447;
      end

       4447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1999] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4448;
      end

       4448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2000] = heapMem[localMem[1982]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4449;
      end

       4449 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2001] = localMem[1929] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4450;
      end

       4450 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2001]) begin
                  heapMem[NArea * localMem[2000] + 0 + i] = heapMem[NArea * localMem[1999] + localMem[1930] + i];
                  updateArrayLength(1, localMem[2000], 0 + i);
                end
              end
              ip = 4451;
      end

       4451 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2002] = heapMem[localMem[1979]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4452;
      end

       4452 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2003] = localMem[2002] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4453;
      end

       4453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2004] = heapMem[localMem[1979]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4454;
      end

       4454 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4455;
      end

       4455 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2005] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4456;
      end

       4456 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4457;
      end

       4457 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2005] >= localMem[2003] ? 4463 : 4458;
      end

       4458 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2006] = heapMem[localMem[2004]*6 + localMem[2005]];
              updateArrayLength(2, 0, 0);
              ip = 4459;
      end

       4459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2006]*6 + 2] = localMem[1979];
              updateArrayLength(1, localMem[2006], 2);
              ip = 4460;
      end

       4460 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4461;
      end

       4461 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2005] = localMem[2005] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4462;
      end

       4462 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4456;
      end

       4463 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4464;
      end

       4464 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2007] = heapMem[localMem[1982]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4465;
      end

       4465 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2008] = localMem[2007] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4466;
      end

       4466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2009] = heapMem[localMem[1982]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4467;
      end

       4467 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4468;
      end

       4468 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2010] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4469;
      end

       4469 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4470;
      end

       4470 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2010] >= localMem[2008] ? 4476 : 4471;
      end

       4471 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2011] = heapMem[localMem[2009]*6 + localMem[2010]];
              updateArrayLength(2, 0, 0);
              ip = 4472;
      end

       4472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2011]*6 + 2] = localMem[1982];
              updateArrayLength(1, localMem[2011], 2);
              ip = 4473;
      end

       4473 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4474;
      end

       4474 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2010] = localMem[2010] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4475;
      end

       4475 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4469;
      end

       4476 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4477;
      end

       4477 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4493;
      end

       4478 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4479;
      end

       4479 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2012] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2012] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2012]] = 0;
              ip = 4480;
      end

       4480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1924]*6 + 6] = localMem[2012];
              updateArrayLength(1, localMem[1924], 6);
              ip = 4481;
      end

       4481 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2013] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4482;
      end

       4482 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2014] = heapMem[localMem[1979]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4483;
      end

       4483 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[2014] + 0 + i] = heapMem[NArea * localMem[2013] + 0 + i];
                  updateArrayLength(1, localMem[2014], 0 + i);
                end
              end
              ip = 4484;
      end

       4484 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2015] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4485;
      end

       4485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2016] = heapMem[localMem[1979]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4486;
      end

       4486 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[2016] + 0 + i] = heapMem[NArea * localMem[2015] + 0 + i];
                  updateArrayLength(1, localMem[2016], 0 + i);
                end
              end
              ip = 4487;
      end

       4487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2017] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4488;
      end

       4488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2018] = heapMem[localMem[1982]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4489;
      end

       4489 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[2018] + 0 + i] = heapMem[NArea * localMem[2017] + localMem[1930] + i];
                  updateArrayLength(1, localMem[2018], 0 + i);
                end
              end
              ip = 4490;
      end

       4490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2019] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4491;
      end

       4491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2020] = heapMem[localMem[1982]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4492;
      end

       4492 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1929]) begin
                  heapMem[NArea * localMem[2020] + 0 + i] = heapMem[NArea * localMem[2019] + localMem[1930] + i];
                  updateArrayLength(1, localMem[2020], 0 + i);
                end
              end
              ip = 4493;
      end

       4493 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4494;
      end

       4494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1979]*6 + 2] = localMem[1924];
              updateArrayLength(1, localMem[1979], 2);
              ip = 4495;
      end

       4495 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1982]*6 + 2] = localMem[1924];
              updateArrayLength(1, localMem[1982], 2);
              ip = 4496;
      end

       4496 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2021] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4497;
      end

       4497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2022] = heapMem[localMem[2021]*6 + localMem[1929]];
              updateArrayLength(2, 0, 0);
              ip = 4498;
      end

       4498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2023] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4499;
      end

       4499 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2024] = heapMem[localMem[2023]*6 + localMem[1929]];
              updateArrayLength(2, 0, 0);
              ip = 4500;
      end

       4500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2025] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4501;
      end

       4501 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2025]*6 + 0] = localMem[2022];
              updateArrayLength(1, localMem[2025], 0);
              ip = 4502;
      end

       4502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2026] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4503;
      end

       4503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2026]*6 + 0] = localMem[2024];
              updateArrayLength(1, localMem[2026], 0);
              ip = 4504;
      end

       4504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2027] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4505;
      end

       4505 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2027]*6 + 0] = localMem[1979];
              updateArrayLength(1, localMem[2027], 0);
              ip = 4506;
      end

       4506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2028] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4507;
      end

       4507 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2028]*6 + 1] = localMem[1982];
              updateArrayLength(1, localMem[2028], 1);
              ip = 4508;
      end

       4508 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1924]*6 + 0] = 1;
              updateArrayLength(1, localMem[1924], 0);
              ip = 4509;
      end

       4509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2029] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4510;
      end

       4510 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2029]] = 1;
              ip = 4511;
      end

       4511 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2030] = heapMem[localMem[1924]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4512;
      end

       4512 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2030]] = 1;
              ip = 4513;
      end

       4513 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2031] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4514;
      end

       4514 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2031]] = 2;
              ip = 4515;
      end

       4515 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4517;
      end

       4516 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4522;
      end

       4517 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4518;
      end

       4518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1925] = 1;
              updateArrayLength(2, 0, 0);
              ip = 4519;
      end

       4519 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4522;
      end

       4520 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4521;
      end

       4521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1925] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4522;
      end

       4522 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4523;
      end

       4523 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4524;
      end

       4524 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4525;
      end

       4525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2032] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4526;
      end

       4526 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4527;
      end

       4527 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2032] >= 99 ? 5025 : 4528;
      end

       4528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2033] = heapMem[localMem[1924]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4529;
      end

       4529 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2034] = localMem[2033] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4530;
      end

       4530 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2035] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4531;
      end

       4531 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2036] = heapMem[localMem[2035]*6 + localMem[2034]];
              updateArrayLength(2, 0, 0);
              ip = 4532;
      end

       4532 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 5 <= localMem[2036] ? 4773 : 4533;
      end

       4533 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2037] = !heapMem[localMem[1924]*6 + 6];
              ip = 4534;
      end

       4534 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2037] == 0 ? 4539 : 4535;
      end

       4535 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 0] = localMem[1924];
              updateArrayLength(1, localMem[1901], 0);
              ip = 4536;
      end

       4536 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 1] = 2;
              updateArrayLength(1, localMem[1901], 1);
              ip = 4537;
      end

       4537 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1901]*6 + 2] = localMem[2033] - 1;
              updateArrayLength(1, localMem[1901], 2);
              ip = 4538;
      end

       4538 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5029;
      end

       4539 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4540;
      end

       4540 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2038] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4541;
      end

       4541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2039] = heapMem[localMem[2038]*6 + localMem[2033]];
              updateArrayLength(2, 0, 0);
              ip = 4542;
      end

       4542 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4543;
      end

       4543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2041] = heapMem[localMem[2039]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4544;
      end

       4544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2042] = heapMem[localMem[2039]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4545;
      end

       4545 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2043] = heapMem[localMem[2042]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4546;
      end

       4546 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2041] <  localMem[2043] ? 4766 : 4547;
      end

       4547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2044] = localMem[2043];
              updateArrayLength(2, 0, 0);
              ip = 4548;
      end

       4548 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2044] = localMem[2044] >> 1;
              ip = 4549;
      end

       4549 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2045] = localMem[2044] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4550;
      end

       4550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2046] = heapMem[localMem[2039]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4551;
      end

       4551 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2046] == 0 ? 4648 : 4552;
      end

       4552 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2047] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2047] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2047]] = 0;
              ip = 4553;
      end

       4553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 0] = localMem[2044];
              updateArrayLength(1, localMem[2047], 0);
              ip = 4554;
      end

       4554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 2] = 0;
              updateArrayLength(1, localMem[2047], 2);
              ip = 4555;
      end

       4555 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2048] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2048] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2048]] = 0;
              ip = 4556;
      end

       4556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 4] = localMem[2048];
              updateArrayLength(1, localMem[2047], 4);
              ip = 4557;
      end

       4557 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2049] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2049] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2049]] = 0;
              ip = 4558;
      end

       4558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 5] = localMem[2049];
              updateArrayLength(1, localMem[2047], 5);
              ip = 4559;
      end

       4559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 6] = 0;
              updateArrayLength(1, localMem[2047], 6);
              ip = 4560;
      end

       4560 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 3] = localMem[2042];
              updateArrayLength(1, localMem[2047], 3);
              ip = 4561;
      end

       4561 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2042]*6 + 1] = heapMem[localMem[2042]*6 + 1] + 1;
              updateArrayLength(1, localMem[2042], 1);
              ip = 4562;
      end

       4562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 1] = heapMem[localMem[2042]*6 + 1];
              updateArrayLength(1, localMem[2047], 1);
              ip = 4563;
      end

       4563 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2050] = !heapMem[localMem[2039]*6 + 6];
              ip = 4564;
      end

       4564 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2050] != 0 ? 4593 : 4565;
      end

       4565 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2051] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2051] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2051]] = 0;
              ip = 4566;
      end

       4566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 6] = localMem[2051];
              updateArrayLength(1, localMem[2047], 6);
              ip = 4567;
      end

       4567 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2052] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4568;
      end

       4568 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2053] = heapMem[localMem[2047]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4569;
      end

       4569 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2053] + 0 + i] = heapMem[NArea * localMem[2052] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2053], 0 + i);
                end
              end
              ip = 4570;
      end

       4570 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2054] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4571;
      end

       4571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2055] = heapMem[localMem[2047]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4572;
      end

       4572 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2055] + 0 + i] = heapMem[NArea * localMem[2054] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2055], 0 + i);
                end
              end
              ip = 4573;
      end

       4573 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2056] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4574;
      end

       4574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2057] = heapMem[localMem[2047]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4575;
      end

       4575 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2058] = localMem[2044] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4576;
      end

       4576 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2058]) begin
                  heapMem[NArea * localMem[2057] + 0 + i] = heapMem[NArea * localMem[2056] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2057], 0 + i);
                end
              end
              ip = 4577;
      end

       4577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2059] = heapMem[localMem[2047]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4578;
      end

       4578 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2060] = localMem[2059] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4579;
      end

       4579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2061] = heapMem[localMem[2047]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4580;
      end

       4580 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4581;
      end

       4581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2062] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4582;
      end

       4582 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4583;
      end

       4583 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2062] >= localMem[2060] ? 4589 : 4584;
      end

       4584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2063] = heapMem[localMem[2061]*6 + localMem[2062]];
              updateArrayLength(2, 0, 0);
              ip = 4585;
      end

       4585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2063]*6 + 2] = localMem[2047];
              updateArrayLength(1, localMem[2063], 2);
              ip = 4586;
      end

       4586 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4587;
      end

       4587 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2062] = localMem[2062] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4588;
      end

       4588 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4582;
      end

       4589 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4590;
      end

       4590 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2064] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4591;
      end

       4591 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2064]] = localMem[2045];
              ip = 4592;
      end

       4592 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4600;
      end

       4593 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4594;
      end

       4594 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2065] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4595;
      end

       4595 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2066] = heapMem[localMem[2047]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4596;
      end

       4596 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2066] + 0 + i] = heapMem[NArea * localMem[2065] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2066], 0 + i);
                end
              end
              ip = 4597;
      end

       4597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2067] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4598;
      end

       4598 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2068] = heapMem[localMem[2047]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4599;
      end

       4599 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2068] + 0 + i] = heapMem[NArea * localMem[2067] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2068], 0 + i);
                end
              end
              ip = 4600;
      end

       4600 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4601;
      end

       4601 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2039]*6 + 0] = localMem[2044];
              updateArrayLength(1, localMem[2039], 0);
              ip = 4602;
      end

       4602 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2047]*6 + 2] = localMem[2046];
              updateArrayLength(1, localMem[2047], 2);
              ip = 4603;
      end

       4603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2069] = heapMem[localMem[2046]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4604;
      end

       4604 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2070] = heapMem[localMem[2046]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4605;
      end

       4605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2071] = heapMem[localMem[2070]*6 + localMem[2069]];
              updateArrayLength(2, 0, 0);
              ip = 4606;
      end

       4606 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2071] != localMem[2039] ? 4625 : 4607;
      end

       4607 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2072] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4608;
      end

       4608 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2073] = heapMem[localMem[2072]*6 + localMem[2044]];
              updateArrayLength(2, 0, 0);
              ip = 4609;
      end

       4609 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2074] = heapMem[localMem[2046]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4610;
      end

       4610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2074]*6 + localMem[2069]] = localMem[2073];
              updateArrayLength(1, localMem[2074], localMem[2069]);
              ip = 4611;
      end

       4611 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2075] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4612;
      end

       4612 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2076] = heapMem[localMem[2075]*6 + localMem[2044]];
              updateArrayLength(2, 0, 0);
              ip = 4613;
      end

       4613 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2077] = heapMem[localMem[2046]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4614;
      end

       4614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2077]*6 + localMem[2069]] = localMem[2076];
              updateArrayLength(1, localMem[2077], localMem[2069]);
              ip = 4615;
      end

       4615 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2078] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4616;
      end

       4616 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2078]] = localMem[2044];
              ip = 4617;
      end

       4617 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2079] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4618;
      end

       4618 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2079]] = localMem[2044];
              ip = 4619;
      end

       4619 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2080] = localMem[2069] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4620;
      end

       4620 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2046]*6 + 0] = localMem[2080];
              updateArrayLength(1, localMem[2046], 0);
              ip = 4621;
      end

       4621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2081] = heapMem[localMem[2046]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4622;
      end

       4622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2081]*6 + localMem[2080]] = localMem[2047];
              updateArrayLength(1, localMem[2081], localMem[2080]);
              ip = 4623;
      end

       4623 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4763;
      end

       4624 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4647;
      end

       4625 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4626;
      end

       4626 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 4627;
      end

       4627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2082] = heapMem[localMem[2046]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4628;
      end

       4628 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2083] = 0; k = arraySizes[localMem[2082]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2082] * NArea + i] == localMem[2039]) localMem[2083] = i + 1;
              end
              ip = 4629;
      end

       4629 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2083] = localMem[2083] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4630;
      end

       4630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2084] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4631;
      end

       4631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2085] = heapMem[localMem[2084]*6 + localMem[2044]];
              updateArrayLength(2, 0, 0);
              ip = 4632;
      end

       4632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2086] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4633;
      end

       4633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2087] = heapMem[localMem[2086]*6 + localMem[2044]];
              updateArrayLength(2, 0, 0);
              ip = 4634;
      end

       4634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2088] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4635;
      end

       4635 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2088]] = localMem[2044];
              ip = 4636;
      end

       4636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2089] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4637;
      end

       4637 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2089]] = localMem[2044];
              ip = 4638;
      end

       4638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2090] = heapMem[localMem[2046]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4639;
      end

       4639 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2090] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2083], localMem[2090], arraySizes[localMem[2090]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2083] && i <= arraySizes[localMem[2090]]) begin
                  heapMem[NArea * localMem[2090] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2090] + localMem[2083]] = localMem[2085];                                    // Insert new value
              arraySizes[localMem[2090]] = arraySizes[localMem[2090]] + 1;                              // Increase array size
              ip = 4640;
      end

       4640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2091] = heapMem[localMem[2046]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4641;
      end

       4641 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2091] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2083], localMem[2091], arraySizes[localMem[2091]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2083] && i <= arraySizes[localMem[2091]]) begin
                  heapMem[NArea * localMem[2091] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2091] + localMem[2083]] = localMem[2087];                                    // Insert new value
              arraySizes[localMem[2091]] = arraySizes[localMem[2091]] + 1;                              // Increase array size
              ip = 4642;
      end

       4642 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2092] = heapMem[localMem[2046]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4643;
      end

       4643 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2093] = localMem[2083] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4644;
      end

       4644 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2092] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2093], localMem[2092], arraySizes[localMem[2092]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2093] && i <= arraySizes[localMem[2092]]) begin
                  heapMem[NArea * localMem[2092] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2092] + localMem[2093]] = localMem[2047];                                    // Insert new value
              arraySizes[localMem[2092]] = arraySizes[localMem[2092]] + 1;                              // Increase array size
              ip = 4645;
      end

       4645 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2046]*6 + 0] = heapMem[localMem[2046]*6 + 0] + 1;
              updateArrayLength(1, localMem[2046], 0);
              ip = 4646;
      end

       4646 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4763;
      end

       4647 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4648;
      end

       4648 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4649;
      end

       4649 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2094] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2094] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2094]] = 0;
              ip = 4650;
      end

       4650 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 0] = localMem[2044];
              updateArrayLength(1, localMem[2094], 0);
              ip = 4651;
      end

       4651 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 2] = 0;
              updateArrayLength(1, localMem[2094], 2);
              ip = 4652;
      end

       4652 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2095] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2095] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2095]] = 0;
              ip = 4653;
      end

       4653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 4] = localMem[2095];
              updateArrayLength(1, localMem[2094], 4);
              ip = 4654;
      end

       4654 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2096] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2096] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2096]] = 0;
              ip = 4655;
      end

       4655 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 5] = localMem[2096];
              updateArrayLength(1, localMem[2094], 5);
              ip = 4656;
      end

       4656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 6] = 0;
              updateArrayLength(1, localMem[2094], 6);
              ip = 4657;
      end

       4657 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 3] = localMem[2042];
              updateArrayLength(1, localMem[2094], 3);
              ip = 4658;
      end

       4658 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2042]*6 + 1] = heapMem[localMem[2042]*6 + 1] + 1;
              updateArrayLength(1, localMem[2042], 1);
              ip = 4659;
      end

       4659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 1] = heapMem[localMem[2042]*6 + 1];
              updateArrayLength(1, localMem[2094], 1);
              ip = 4660;
      end

       4660 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2097] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2097] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2097]] = 0;
              ip = 4661;
      end

       4661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 0] = localMem[2044];
              updateArrayLength(1, localMem[2097], 0);
              ip = 4662;
      end

       4662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 2] = 0;
              updateArrayLength(1, localMem[2097], 2);
              ip = 4663;
      end

       4663 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2098] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2098] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2098]] = 0;
              ip = 4664;
      end

       4664 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 4] = localMem[2098];
              updateArrayLength(1, localMem[2097], 4);
              ip = 4665;
      end

       4665 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2099] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2099] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2099]] = 0;
              ip = 4666;
      end

       4666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 5] = localMem[2099];
              updateArrayLength(1, localMem[2097], 5);
              ip = 4667;
      end

       4667 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 6] = 0;
              updateArrayLength(1, localMem[2097], 6);
              ip = 4668;
      end

       4668 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 3] = localMem[2042];
              updateArrayLength(1, localMem[2097], 3);
              ip = 4669;
      end

       4669 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2042]*6 + 1] = heapMem[localMem[2042]*6 + 1] + 1;
              updateArrayLength(1, localMem[2042], 1);
              ip = 4670;
      end

       4670 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 1] = heapMem[localMem[2042]*6 + 1];
              updateArrayLength(1, localMem[2097], 1);
              ip = 4671;
      end

       4671 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2100] = !heapMem[localMem[2039]*6 + 6];
              ip = 4672;
      end

       4672 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2100] != 0 ? 4724 : 4673;
      end

       4673 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2101] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2101] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2101]] = 0;
              ip = 4674;
      end

       4674 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 6] = localMem[2101];
              updateArrayLength(1, localMem[2094], 6);
              ip = 4675;
      end

       4675 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2102] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2102] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2102]] = 0;
              ip = 4676;
      end

       4676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 6] = localMem[2102];
              updateArrayLength(1, localMem[2097], 6);
              ip = 4677;
      end

       4677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2103] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4678;
      end

       4678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2104] = heapMem[localMem[2094]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4679;
      end

       4679 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2104] + 0 + i] = heapMem[NArea * localMem[2103] + 0 + i];
                  updateArrayLength(1, localMem[2104], 0 + i);
                end
              end
              ip = 4680;
      end

       4680 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2105] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4681;
      end

       4681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2106] = heapMem[localMem[2094]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4682;
      end

       4682 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2106] + 0 + i] = heapMem[NArea * localMem[2105] + 0 + i];
                  updateArrayLength(1, localMem[2106], 0 + i);
                end
              end
              ip = 4683;
      end

       4683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2107] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4684;
      end

       4684 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2108] = heapMem[localMem[2094]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4685;
      end

       4685 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2109] = localMem[2044] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4686;
      end

       4686 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2109]) begin
                  heapMem[NArea * localMem[2108] + 0 + i] = heapMem[NArea * localMem[2107] + 0 + i];
                  updateArrayLength(1, localMem[2108], 0 + i);
                end
              end
              ip = 4687;
      end

       4687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2110] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4688;
      end

       4688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2111] = heapMem[localMem[2097]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4689;
      end

       4689 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2111] + 0 + i] = heapMem[NArea * localMem[2110] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2111], 0 + i);
                end
              end
              ip = 4690;
      end

       4690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2112] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4691;
      end

       4691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2113] = heapMem[localMem[2097]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4692;
      end

       4692 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2113] + 0 + i] = heapMem[NArea * localMem[2112] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2113], 0 + i);
                end
              end
              ip = 4693;
      end

       4693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2114] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4694;
      end

       4694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2115] = heapMem[localMem[2097]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4695;
      end

       4695 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2116] = localMem[2044] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4696;
      end

       4696 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2116]) begin
                  heapMem[NArea * localMem[2115] + 0 + i] = heapMem[NArea * localMem[2114] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2115], 0 + i);
                end
              end
              ip = 4697;
      end

       4697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2117] = heapMem[localMem[2094]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4698;
      end

       4698 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2118] = localMem[2117] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4699;
      end

       4699 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2119] = heapMem[localMem[2094]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4700;
      end

       4700 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4701;
      end

       4701 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2120] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4702;
      end

       4702 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4703;
      end

       4703 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2120] >= localMem[2118] ? 4709 : 4704;
      end

       4704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2121] = heapMem[localMem[2119]*6 + localMem[2120]];
              updateArrayLength(2, 0, 0);
              ip = 4705;
      end

       4705 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2121]*6 + 2] = localMem[2094];
              updateArrayLength(1, localMem[2121], 2);
              ip = 4706;
      end

       4706 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4707;
      end

       4707 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2120] = localMem[2120] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4708;
      end

       4708 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4702;
      end

       4709 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4710;
      end

       4710 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2122] = heapMem[localMem[2097]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4711;
      end

       4711 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2123] = localMem[2122] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4712;
      end

       4712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2124] = heapMem[localMem[2097]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4713;
      end

       4713 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4714;
      end

       4714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2125] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4715;
      end

       4715 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4716;
      end

       4716 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2125] >= localMem[2123] ? 4722 : 4717;
      end

       4717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2126] = heapMem[localMem[2124]*6 + localMem[2125]];
              updateArrayLength(2, 0, 0);
              ip = 4718;
      end

       4718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2126]*6 + 2] = localMem[2097];
              updateArrayLength(1, localMem[2126], 2);
              ip = 4719;
      end

       4719 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4720;
      end

       4720 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2125] = localMem[2125] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4721;
      end

       4721 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4715;
      end

       4722 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4723;
      end

       4723 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4739;
      end

       4724 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4725;
      end

       4725 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2127] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2127] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2127]] = 0;
              ip = 4726;
      end

       4726 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2039]*6 + 6] = localMem[2127];
              updateArrayLength(1, localMem[2039], 6);
              ip = 4727;
      end

       4727 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2128] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4728;
      end

       4728 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2129] = heapMem[localMem[2094]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4729;
      end

       4729 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2129] + 0 + i] = heapMem[NArea * localMem[2128] + 0 + i];
                  updateArrayLength(1, localMem[2129], 0 + i);
                end
              end
              ip = 4730;
      end

       4730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2130] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4731;
      end

       4731 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2131] = heapMem[localMem[2094]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4732;
      end

       4732 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2131] + 0 + i] = heapMem[NArea * localMem[2130] + 0 + i];
                  updateArrayLength(1, localMem[2131], 0 + i);
                end
              end
              ip = 4733;
      end

       4733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2132] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4734;
      end

       4734 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2133] = heapMem[localMem[2097]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4735;
      end

       4735 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2133] + 0 + i] = heapMem[NArea * localMem[2132] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2133], 0 + i);
                end
              end
              ip = 4736;
      end

       4736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2134] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4737;
      end

       4737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2135] = heapMem[localMem[2097]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4738;
      end

       4738 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2044]) begin
                  heapMem[NArea * localMem[2135] + 0 + i] = heapMem[NArea * localMem[2134] + localMem[2045] + i];
                  updateArrayLength(1, localMem[2135], 0 + i);
                end
              end
              ip = 4739;
      end

       4739 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4740;
      end

       4740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2094]*6 + 2] = localMem[2039];
              updateArrayLength(1, localMem[2094], 2);
              ip = 4741;
      end

       4741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2097]*6 + 2] = localMem[2039];
              updateArrayLength(1, localMem[2097], 2);
              ip = 4742;
      end

       4742 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2136] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4743;
      end

       4743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2137] = heapMem[localMem[2136]*6 + localMem[2044]];
              updateArrayLength(2, 0, 0);
              ip = 4744;
      end

       4744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2138] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4745;
      end

       4745 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2139] = heapMem[localMem[2138]*6 + localMem[2044]];
              updateArrayLength(2, 0, 0);
              ip = 4746;
      end

       4746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2140] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4747;
      end

       4747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2140]*6 + 0] = localMem[2137];
              updateArrayLength(1, localMem[2140], 0);
              ip = 4748;
      end

       4748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2141] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4749;
      end

       4749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2141]*6 + 0] = localMem[2139];
              updateArrayLength(1, localMem[2141], 0);
              ip = 4750;
      end

       4750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2142] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4751;
      end

       4751 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2142]*6 + 0] = localMem[2094];
              updateArrayLength(1, localMem[2142], 0);
              ip = 4752;
      end

       4752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2143] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4753;
      end

       4753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2143]*6 + 1] = localMem[2097];
              updateArrayLength(1, localMem[2143], 1);
              ip = 4754;
      end

       4754 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2039]*6 + 0] = 1;
              updateArrayLength(1, localMem[2039], 0);
              ip = 4755;
      end

       4755 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2144] = heapMem[localMem[2039]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4756;
      end

       4756 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2144]] = 1;
              ip = 4757;
      end

       4757 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2145] = heapMem[localMem[2039]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4758;
      end

       4758 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2145]] = 1;
              ip = 4759;
      end

       4759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2146] = heapMem[localMem[2039]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4760;
      end

       4760 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2146]] = 2;
              ip = 4761;
      end

       4761 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4763;
      end

       4762 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4768;
      end

       4763 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4764;
      end

       4764 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2040] = 1;
              updateArrayLength(2, 0, 0);
              ip = 4765;
      end

       4765 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4768;
      end

       4766 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4767;
      end

       4767 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2040] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4768;
      end

       4768 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4769;
      end

       4769 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2040] != 0 ? 4771 : 4770;
      end

       4770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1924] = localMem[2039];
              updateArrayLength(2, 0, 0);
              ip = 4771;
      end

       4771 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4772;
      end

       4772 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5022;
      end

       4773 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4774;
      end

       4774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2147] = heapMem[localMem[1924]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4775;
      end

       4775 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2148] = 0; k = arraySizes[localMem[2147]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2147] * NArea + i] == 5) localMem[2148] = i + 1;
              end
              ip = 4776;
      end

       4776 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2148] == 0 ? 4781 : 4777;
      end

       4777 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 0] = localMem[1924];
              updateArrayLength(1, localMem[1901], 0);
              ip = 4778;
      end

       4778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 1] = 1;
              updateArrayLength(1, localMem[1901], 1);
              ip = 4779;
      end

       4779 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1901]*6 + 2] = localMem[2148] - 1;
              updateArrayLength(1, localMem[1901], 2);
              ip = 4780;
      end

       4780 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5029;
      end

       4781 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4782;
      end

       4782 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[2147]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2147] * NArea + i] < 5) j = j + 1;
              end
              localMem[2149] = j;
              ip = 4783;
      end

       4783 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2150] = !heapMem[localMem[1924]*6 + 6];
              ip = 4784;
      end

       4784 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2150] == 0 ? 4789 : 4785;
      end

       4785 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 0] = localMem[1924];
              updateArrayLength(1, localMem[1901], 0);
              ip = 4786;
      end

       4786 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 1] = 0;
              updateArrayLength(1, localMem[1901], 1);
              ip = 4787;
      end

       4787 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*6 + 2] = localMem[2149];
              updateArrayLength(1, localMem[1901], 2);
              ip = 4788;
      end

       4788 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5029;
      end

       4789 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4790;
      end

       4790 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2151] = heapMem[localMem[1924]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4791;
      end

       4791 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2152] = heapMem[localMem[2151]*6 + localMem[2149]];
              updateArrayLength(2, 0, 0);
              ip = 4792;
      end

       4792 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4793;
      end

       4793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2154] = heapMem[localMem[2152]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4794;
      end

       4794 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2155] = heapMem[localMem[2152]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4795;
      end

       4795 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2156] = heapMem[localMem[2155]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4796;
      end

       4796 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2154] <  localMem[2156] ? 5016 : 4797;
      end

       4797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2157] = localMem[2156];
              updateArrayLength(2, 0, 0);
              ip = 4798;
      end

       4798 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2157] = localMem[2157] >> 1;
              ip = 4799;
      end

       4799 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2158] = localMem[2157] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4800;
      end

       4800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2159] = heapMem[localMem[2152]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4801;
      end

       4801 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2159] == 0 ? 4898 : 4802;
      end

       4802 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2160] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2160] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2160]] = 0;
              ip = 4803;
      end

       4803 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 0] = localMem[2157];
              updateArrayLength(1, localMem[2160], 0);
              ip = 4804;
      end

       4804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 2] = 0;
              updateArrayLength(1, localMem[2160], 2);
              ip = 4805;
      end

       4805 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2161] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2161] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2161]] = 0;
              ip = 4806;
      end

       4806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 4] = localMem[2161];
              updateArrayLength(1, localMem[2160], 4);
              ip = 4807;
      end

       4807 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2162] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2162] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2162]] = 0;
              ip = 4808;
      end

       4808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 5] = localMem[2162];
              updateArrayLength(1, localMem[2160], 5);
              ip = 4809;
      end

       4809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 6] = 0;
              updateArrayLength(1, localMem[2160], 6);
              ip = 4810;
      end

       4810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 3] = localMem[2155];
              updateArrayLength(1, localMem[2160], 3);
              ip = 4811;
      end

       4811 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2155]*6 + 1] = heapMem[localMem[2155]*6 + 1] + 1;
              updateArrayLength(1, localMem[2155], 1);
              ip = 4812;
      end

       4812 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 1] = heapMem[localMem[2155]*6 + 1];
              updateArrayLength(1, localMem[2160], 1);
              ip = 4813;
      end

       4813 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2163] = !heapMem[localMem[2152]*6 + 6];
              ip = 4814;
      end

       4814 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2163] != 0 ? 4843 : 4815;
      end

       4815 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2164] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2164] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2164]] = 0;
              ip = 4816;
      end

       4816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 6] = localMem[2164];
              updateArrayLength(1, localMem[2160], 6);
              ip = 4817;
      end

       4817 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2165] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4818;
      end

       4818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2166] = heapMem[localMem[2160]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4819;
      end

       4819 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2166] + 0 + i] = heapMem[NArea * localMem[2165] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2166], 0 + i);
                end
              end
              ip = 4820;
      end

       4820 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2167] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4821;
      end

       4821 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2168] = heapMem[localMem[2160]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4822;
      end

       4822 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2168] + 0 + i] = heapMem[NArea * localMem[2167] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2168], 0 + i);
                end
              end
              ip = 4823;
      end

       4823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2169] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4824;
      end

       4824 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2170] = heapMem[localMem[2160]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4825;
      end

       4825 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2171] = localMem[2157] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4826;
      end

       4826 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2171]) begin
                  heapMem[NArea * localMem[2170] + 0 + i] = heapMem[NArea * localMem[2169] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2170], 0 + i);
                end
              end
              ip = 4827;
      end

       4827 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2172] = heapMem[localMem[2160]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4828;
      end

       4828 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2173] = localMem[2172] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4829;
      end

       4829 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2174] = heapMem[localMem[2160]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4830;
      end

       4830 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4831;
      end

       4831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2175] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4832;
      end

       4832 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4833;
      end

       4833 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2175] >= localMem[2173] ? 4839 : 4834;
      end

       4834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2176] = heapMem[localMem[2174]*6 + localMem[2175]];
              updateArrayLength(2, 0, 0);
              ip = 4835;
      end

       4835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2176]*6 + 2] = localMem[2160];
              updateArrayLength(1, localMem[2176], 2);
              ip = 4836;
      end

       4836 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4837;
      end

       4837 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2175] = localMem[2175] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4838;
      end

       4838 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4832;
      end

       4839 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4840;
      end

       4840 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2177] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4841;
      end

       4841 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2177]] = localMem[2158];
              ip = 4842;
      end

       4842 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4850;
      end

       4843 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4844;
      end

       4844 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2178] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4845;
      end

       4845 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2179] = heapMem[localMem[2160]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4846;
      end

       4846 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2179] + 0 + i] = heapMem[NArea * localMem[2178] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2179], 0 + i);
                end
              end
              ip = 4847;
      end

       4847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2180] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4848;
      end

       4848 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2181] = heapMem[localMem[2160]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4849;
      end

       4849 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2181] + 0 + i] = heapMem[NArea * localMem[2180] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2181], 0 + i);
                end
              end
              ip = 4850;
      end

       4850 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4851;
      end

       4851 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2152]*6 + 0] = localMem[2157];
              updateArrayLength(1, localMem[2152], 0);
              ip = 4852;
      end

       4852 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2160]*6 + 2] = localMem[2159];
              updateArrayLength(1, localMem[2160], 2);
              ip = 4853;
      end

       4853 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2182] = heapMem[localMem[2159]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4854;
      end

       4854 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2183] = heapMem[localMem[2159]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4855;
      end

       4855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2184] = heapMem[localMem[2183]*6 + localMem[2182]];
              updateArrayLength(2, 0, 0);
              ip = 4856;
      end

       4856 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2184] != localMem[2152] ? 4875 : 4857;
      end

       4857 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2185] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4858;
      end

       4858 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2186] = heapMem[localMem[2185]*6 + localMem[2157]];
              updateArrayLength(2, 0, 0);
              ip = 4859;
      end

       4859 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2187] = heapMem[localMem[2159]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4860;
      end

       4860 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2187]*6 + localMem[2182]] = localMem[2186];
              updateArrayLength(1, localMem[2187], localMem[2182]);
              ip = 4861;
      end

       4861 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2188] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4862;
      end

       4862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2189] = heapMem[localMem[2188]*6 + localMem[2157]];
              updateArrayLength(2, 0, 0);
              ip = 4863;
      end

       4863 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2190] = heapMem[localMem[2159]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4864;
      end

       4864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2190]*6 + localMem[2182]] = localMem[2189];
              updateArrayLength(1, localMem[2190], localMem[2182]);
              ip = 4865;
      end

       4865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2191] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4866;
      end

       4866 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2191]] = localMem[2157];
              ip = 4867;
      end

       4867 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2192] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4868;
      end

       4868 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2192]] = localMem[2157];
              ip = 4869;
      end

       4869 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2193] = localMem[2182] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4870;
      end

       4870 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2159]*6 + 0] = localMem[2193];
              updateArrayLength(1, localMem[2159], 0);
              ip = 4871;
      end

       4871 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2194] = heapMem[localMem[2159]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4872;
      end

       4872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2194]*6 + localMem[2193]] = localMem[2160];
              updateArrayLength(1, localMem[2194], localMem[2193]);
              ip = 4873;
      end

       4873 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5013;
      end

       4874 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4897;
      end

       4875 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4876;
      end

       4876 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 4877;
      end

       4877 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2195] = heapMem[localMem[2159]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4878;
      end

       4878 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2196] = 0; k = arraySizes[localMem[2195]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2195] * NArea + i] == localMem[2152]) localMem[2196] = i + 1;
              end
              ip = 4879;
      end

       4879 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2196] = localMem[2196] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4880;
      end

       4880 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2197] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4881;
      end

       4881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2198] = heapMem[localMem[2197]*6 + localMem[2157]];
              updateArrayLength(2, 0, 0);
              ip = 4882;
      end

       4882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2199] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4883;
      end

       4883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2200] = heapMem[localMem[2199]*6 + localMem[2157]];
              updateArrayLength(2, 0, 0);
              ip = 4884;
      end

       4884 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2201] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4885;
      end

       4885 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2201]] = localMem[2157];
              ip = 4886;
      end

       4886 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2202] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4887;
      end

       4887 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2202]] = localMem[2157];
              ip = 4888;
      end

       4888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2203] = heapMem[localMem[2159]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4889;
      end

       4889 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2203] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2196], localMem[2203], arraySizes[localMem[2203]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2196] && i <= arraySizes[localMem[2203]]) begin
                  heapMem[NArea * localMem[2203] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2203] + localMem[2196]] = localMem[2198];                                    // Insert new value
              arraySizes[localMem[2203]] = arraySizes[localMem[2203]] + 1;                              // Increase array size
              ip = 4890;
      end

       4890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2204] = heapMem[localMem[2159]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4891;
      end

       4891 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2204] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2196], localMem[2204], arraySizes[localMem[2204]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2196] && i <= arraySizes[localMem[2204]]) begin
                  heapMem[NArea * localMem[2204] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2204] + localMem[2196]] = localMem[2200];                                    // Insert new value
              arraySizes[localMem[2204]] = arraySizes[localMem[2204]] + 1;                              // Increase array size
              ip = 4892;
      end

       4892 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2205] = heapMem[localMem[2159]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4893;
      end

       4893 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2206] = localMem[2196] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4894;
      end

       4894 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2205] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2206], localMem[2205], arraySizes[localMem[2205]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2206] && i <= arraySizes[localMem[2205]]) begin
                  heapMem[NArea * localMem[2205] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2205] + localMem[2206]] = localMem[2160];                                    // Insert new value
              arraySizes[localMem[2205]] = arraySizes[localMem[2205]] + 1;                              // Increase array size
              ip = 4895;
      end

       4895 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2159]*6 + 0] = heapMem[localMem[2159]*6 + 0] + 1;
              updateArrayLength(1, localMem[2159], 0);
              ip = 4896;
      end

       4896 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5013;
      end

       4897 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4898;
      end

       4898 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4899;
      end

       4899 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2207] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2207] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2207]] = 0;
              ip = 4900;
      end

       4900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 0] = localMem[2157];
              updateArrayLength(1, localMem[2207], 0);
              ip = 4901;
      end

       4901 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 2] = 0;
              updateArrayLength(1, localMem[2207], 2);
              ip = 4902;
      end

       4902 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2208] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2208] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2208]] = 0;
              ip = 4903;
      end

       4903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 4] = localMem[2208];
              updateArrayLength(1, localMem[2207], 4);
              ip = 4904;
      end

       4904 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2209] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2209] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2209]] = 0;
              ip = 4905;
      end

       4905 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 5] = localMem[2209];
              updateArrayLength(1, localMem[2207], 5);
              ip = 4906;
      end

       4906 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 6] = 0;
              updateArrayLength(1, localMem[2207], 6);
              ip = 4907;
      end

       4907 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 3] = localMem[2155];
              updateArrayLength(1, localMem[2207], 3);
              ip = 4908;
      end

       4908 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2155]*6 + 1] = heapMem[localMem[2155]*6 + 1] + 1;
              updateArrayLength(1, localMem[2155], 1);
              ip = 4909;
      end

       4909 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 1] = heapMem[localMem[2155]*6 + 1];
              updateArrayLength(1, localMem[2207], 1);
              ip = 4910;
      end

       4910 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2210] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2210] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2210]] = 0;
              ip = 4911;
      end

       4911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 0] = localMem[2157];
              updateArrayLength(1, localMem[2210], 0);
              ip = 4912;
      end

       4912 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 2] = 0;
              updateArrayLength(1, localMem[2210], 2);
              ip = 4913;
      end

       4913 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2211] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2211] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2211]] = 0;
              ip = 4914;
      end

       4914 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 4] = localMem[2211];
              updateArrayLength(1, localMem[2210], 4);
              ip = 4915;
      end

       4915 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2212] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2212] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2212]] = 0;
              ip = 4916;
      end

       4916 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 5] = localMem[2212];
              updateArrayLength(1, localMem[2210], 5);
              ip = 4917;
      end

       4917 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 6] = 0;
              updateArrayLength(1, localMem[2210], 6);
              ip = 4918;
      end

       4918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 3] = localMem[2155];
              updateArrayLength(1, localMem[2210], 3);
              ip = 4919;
      end

       4919 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2155]*6 + 1] = heapMem[localMem[2155]*6 + 1] + 1;
              updateArrayLength(1, localMem[2155], 1);
              ip = 4920;
      end

       4920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 1] = heapMem[localMem[2155]*6 + 1];
              updateArrayLength(1, localMem[2210], 1);
              ip = 4921;
      end

       4921 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2213] = !heapMem[localMem[2152]*6 + 6];
              ip = 4922;
      end

       4922 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2213] != 0 ? 4974 : 4923;
      end

       4923 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2214] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2214] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2214]] = 0;
              ip = 4924;
      end

       4924 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 6] = localMem[2214];
              updateArrayLength(1, localMem[2207], 6);
              ip = 4925;
      end

       4925 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2215] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2215] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2215]] = 0;
              ip = 4926;
      end

       4926 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 6] = localMem[2215];
              updateArrayLength(1, localMem[2210], 6);
              ip = 4927;
      end

       4927 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2216] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4928;
      end

       4928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2217] = heapMem[localMem[2207]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4929;
      end

       4929 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2217] + 0 + i] = heapMem[NArea * localMem[2216] + 0 + i];
                  updateArrayLength(1, localMem[2217], 0 + i);
                end
              end
              ip = 4930;
      end

       4930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2218] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4931;
      end

       4931 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2219] = heapMem[localMem[2207]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4932;
      end

       4932 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2219] + 0 + i] = heapMem[NArea * localMem[2218] + 0 + i];
                  updateArrayLength(1, localMem[2219], 0 + i);
                end
              end
              ip = 4933;
      end

       4933 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2220] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4934;
      end

       4934 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2221] = heapMem[localMem[2207]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4935;
      end

       4935 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2222] = localMem[2157] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4936;
      end

       4936 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2222]) begin
                  heapMem[NArea * localMem[2221] + 0 + i] = heapMem[NArea * localMem[2220] + 0 + i];
                  updateArrayLength(1, localMem[2221], 0 + i);
                end
              end
              ip = 4937;
      end

       4937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2223] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4938;
      end

       4938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2224] = heapMem[localMem[2210]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4939;
      end

       4939 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2224] + 0 + i] = heapMem[NArea * localMem[2223] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2224], 0 + i);
                end
              end
              ip = 4940;
      end

       4940 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2225] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4941;
      end

       4941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2226] = heapMem[localMem[2210]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4942;
      end

       4942 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2226] + 0 + i] = heapMem[NArea * localMem[2225] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2226], 0 + i);
                end
              end
              ip = 4943;
      end

       4943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2227] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4944;
      end

       4944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2228] = heapMem[localMem[2210]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4945;
      end

       4945 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2229] = localMem[2157] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4946;
      end

       4946 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2229]) begin
                  heapMem[NArea * localMem[2228] + 0 + i] = heapMem[NArea * localMem[2227] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2228], 0 + i);
                end
              end
              ip = 4947;
      end

       4947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2230] = heapMem[localMem[2207]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4948;
      end

       4948 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2231] = localMem[2230] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4949;
      end

       4949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2232] = heapMem[localMem[2207]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4950;
      end

       4950 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4951;
      end

       4951 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2233] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4952;
      end

       4952 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4953;
      end

       4953 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2233] >= localMem[2231] ? 4959 : 4954;
      end

       4954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2234] = heapMem[localMem[2232]*6 + localMem[2233]];
              updateArrayLength(2, 0, 0);
              ip = 4955;
      end

       4955 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2234]*6 + 2] = localMem[2207];
              updateArrayLength(1, localMem[2234], 2);
              ip = 4956;
      end

       4956 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4957;
      end

       4957 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2233] = localMem[2233] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4958;
      end

       4958 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4952;
      end

       4959 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4960;
      end

       4960 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2235] = heapMem[localMem[2210]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4961;
      end

       4961 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2236] = localMem[2235] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4962;
      end

       4962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2237] = heapMem[localMem[2210]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4963;
      end

       4963 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4964;
      end

       4964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2238] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4965;
      end

       4965 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4966;
      end

       4966 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2238] >= localMem[2236] ? 4972 : 4967;
      end

       4967 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2239] = heapMem[localMem[2237]*6 + localMem[2238]];
              updateArrayLength(2, 0, 0);
              ip = 4968;
      end

       4968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2239]*6 + 2] = localMem[2210];
              updateArrayLength(1, localMem[2239], 2);
              ip = 4969;
      end

       4969 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4970;
      end

       4970 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2238] = localMem[2238] + 1;
              updateArrayLength(2, 0, 0);
              ip = 4971;
      end

       4971 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4965;
      end

       4972 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4973;
      end

       4973 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4989;
      end

       4974 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4975;
      end

       4975 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2240] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2240] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2240]] = 0;
              ip = 4976;
      end

       4976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2152]*6 + 6] = localMem[2240];
              updateArrayLength(1, localMem[2152], 6);
              ip = 4977;
      end

       4977 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2241] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4978;
      end

       4978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2242] = heapMem[localMem[2207]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4979;
      end

       4979 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2242] + 0 + i] = heapMem[NArea * localMem[2241] + 0 + i];
                  updateArrayLength(1, localMem[2242], 0 + i);
                end
              end
              ip = 4980;
      end

       4980 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2243] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4981;
      end

       4981 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2244] = heapMem[localMem[2207]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4982;
      end

       4982 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2244] + 0 + i] = heapMem[NArea * localMem[2243] + 0 + i];
                  updateArrayLength(1, localMem[2244], 0 + i);
                end
              end
              ip = 4983;
      end

       4983 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2245] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4984;
      end

       4984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2246] = heapMem[localMem[2210]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4985;
      end

       4985 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2246] + 0 + i] = heapMem[NArea * localMem[2245] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2246], 0 + i);
                end
              end
              ip = 4986;
      end

       4986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2247] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4987;
      end

       4987 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2248] = heapMem[localMem[2210]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4988;
      end

       4988 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2157]) begin
                  heapMem[NArea * localMem[2248] + 0 + i] = heapMem[NArea * localMem[2247] + localMem[2158] + i];
                  updateArrayLength(1, localMem[2248], 0 + i);
                end
              end
              ip = 4989;
      end

       4989 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4990;
      end

       4990 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2207]*6 + 2] = localMem[2152];
              updateArrayLength(1, localMem[2207], 2);
              ip = 4991;
      end

       4991 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2210]*6 + 2] = localMem[2152];
              updateArrayLength(1, localMem[2210], 2);
              ip = 4992;
      end

       4992 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2249] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4993;
      end

       4993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2250] = heapMem[localMem[2249]*6 + localMem[2157]];
              updateArrayLength(2, 0, 0);
              ip = 4994;
      end

       4994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2251] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4995;
      end

       4995 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2252] = heapMem[localMem[2251]*6 + localMem[2157]];
              updateArrayLength(2, 0, 0);
              ip = 4996;
      end

       4996 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2253] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4997;
      end

       4997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2253]*6 + 0] = localMem[2250];
              updateArrayLength(1, localMem[2253], 0);
              ip = 4998;
      end

       4998 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2254] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 4999;
      end

       4999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2254]*6 + 0] = localMem[2252];
              updateArrayLength(1, localMem[2254], 0);
              ip = 5000;
      end

       5000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2255] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5001;
      end

       5001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2255]*6 + 0] = localMem[2207];
              updateArrayLength(1, localMem[2255], 0);
              ip = 5002;
      end

       5002 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2256] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5003;
      end

       5003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2256]*6 + 1] = localMem[2210];
              updateArrayLength(1, localMem[2256], 1);
              ip = 5004;
      end

       5004 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2152]*6 + 0] = 1;
              updateArrayLength(1, localMem[2152], 0);
              ip = 5005;
      end

       5005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2257] = heapMem[localMem[2152]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5006;
      end

       5006 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2257]] = 1;
              ip = 5007;
      end

       5007 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2258] = heapMem[localMem[2152]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5008;
      end

       5008 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2258]] = 1;
              ip = 5009;
      end

       5009 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2259] = heapMem[localMem[2152]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5010;
      end

       5010 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2259]] = 2;
              ip = 5011;
      end

       5011 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5013;
      end

       5012 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5018;
      end

       5013 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5014;
      end

       5014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2153] = 1;
              updateArrayLength(2, 0, 0);
              ip = 5015;
      end

       5015 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5018;
      end

       5016 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5017;
      end

       5017 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2153] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5018;
      end

       5018 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5019;
      end

       5019 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2153] != 0 ? 5021 : 5020;
      end

       5020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1924] = localMem[2152];
              updateArrayLength(2, 0, 0);
              ip = 5021;
      end

       5021 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5022;
      end

       5022 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5023;
      end

       5023 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2032] = localMem[2032] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5024;
      end

       5024 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4526;
      end

       5025 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5026;
      end

       5026 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
            ip = 5027;
      end

       5027 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5028;
      end

       5028 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5029;
      end

       5029 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5030;
      end

       5030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2260] = heapMem[localMem[1901]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5031;
      end

       5031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2261] = heapMem[localMem[1901]*6 + 1];
              updateArrayLength(2, 0, 0);
              ip = 5032;
      end

       5032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2262] = heapMem[localMem[1901]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5033;
      end

       5033 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2261] != 1 ? 5037 : 5034;
      end

       5034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2263] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5035;
      end

       5035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2263]*6 + localMem[2262]] = 55;
              updateArrayLength(1, localMem[2263], localMem[2262]);
              ip = 5036;
      end

       5036 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5283;
      end

       5037 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5038;
      end

       5038 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2261] != 2 ? 5046 : 5039;
      end

       5039 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2264] = localMem[2262] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5040;
      end

       5040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2265] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5041;
      end

       5041 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2265] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2264], localMem[2265], arraySizes[localMem[2265]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2264] && i <= arraySizes[localMem[2265]]) begin
                  heapMem[NArea * localMem[2265] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2265] + localMem[2264]] = 5;                                    // Insert new value
              arraySizes[localMem[2265]] = arraySizes[localMem[2265]] + 1;                              // Increase array size
              ip = 5042;
      end

       5042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2266] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5043;
      end

       5043 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2266] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2264], localMem[2266], arraySizes[localMem[2266]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2264] && i <= arraySizes[localMem[2266]]) begin
                  heapMem[NArea * localMem[2266] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2266] + localMem[2264]] = 55;                                    // Insert new value
              arraySizes[localMem[2266]] = arraySizes[localMem[2266]] + 1;                              // Increase array size
              ip = 5044;
      end

       5044 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2260]*6 + 0] = heapMem[localMem[2260]*6 + 0] + 1;
              updateArrayLength(1, localMem[2260], 0);
              ip = 5045;
      end

       5045 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5052;
      end

       5046 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5047;
      end

       5047 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2267] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5048;
      end

       5048 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2267] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2262], localMem[2267], arraySizes[localMem[2267]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2262] && i <= arraySizes[localMem[2267]]) begin
                  heapMem[NArea * localMem[2267] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2267] + localMem[2262]] = 5;                                    // Insert new value
              arraySizes[localMem[2267]] = arraySizes[localMem[2267]] + 1;                              // Increase array size
              ip = 5049;
      end

       5049 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2268] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5050;
      end

       5050 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2268] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2262], localMem[2268], arraySizes[localMem[2268]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2262] && i <= arraySizes[localMem[2268]]) begin
                  heapMem[NArea * localMem[2268] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2268] + localMem[2262]] = 55;                                    // Insert new value
              arraySizes[localMem[2268]] = arraySizes[localMem[2268]] + 1;                              // Increase array size
              ip = 5051;
      end

       5051 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2260]*6 + 0] = heapMem[localMem[2260]*6 + 0] + 1;
              updateArrayLength(1, localMem[2260], 0);
              ip = 5052;
      end

       5052 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5053;
      end

       5053 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 5054;
      end

       5054 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5055;
      end

       5055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2270] = heapMem[localMem[2260]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5056;
      end

       5056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2271] = heapMem[localMem[2260]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5057;
      end

       5057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2272] = heapMem[localMem[2271]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5058;
      end

       5058 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2270] <  localMem[2272] ? 5278 : 5059;
      end

       5059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2273] = localMem[2272];
              updateArrayLength(2, 0, 0);
              ip = 5060;
      end

       5060 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2273] = localMem[2273] >> 1;
              ip = 5061;
      end

       5061 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2274] = localMem[2273] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5062;
      end

       5062 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2275] = heapMem[localMem[2260]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5063;
      end

       5063 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2275] == 0 ? 5160 : 5064;
      end

       5064 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2276] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2276] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2276]] = 0;
              ip = 5065;
      end

       5065 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 0] = localMem[2273];
              updateArrayLength(1, localMem[2276], 0);
              ip = 5066;
      end

       5066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 2] = 0;
              updateArrayLength(1, localMem[2276], 2);
              ip = 5067;
      end

       5067 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2277] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2277] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2277]] = 0;
              ip = 5068;
      end

       5068 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 4] = localMem[2277];
              updateArrayLength(1, localMem[2276], 4);
              ip = 5069;
      end

       5069 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2278] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2278] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2278]] = 0;
              ip = 5070;
      end

       5070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 5] = localMem[2278];
              updateArrayLength(1, localMem[2276], 5);
              ip = 5071;
      end

       5071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 6] = 0;
              updateArrayLength(1, localMem[2276], 6);
              ip = 5072;
      end

       5072 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 3] = localMem[2271];
              updateArrayLength(1, localMem[2276], 3);
              ip = 5073;
      end

       5073 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2271]*6 + 1] = heapMem[localMem[2271]*6 + 1] + 1;
              updateArrayLength(1, localMem[2271], 1);
              ip = 5074;
      end

       5074 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 1] = heapMem[localMem[2271]*6 + 1];
              updateArrayLength(1, localMem[2276], 1);
              ip = 5075;
      end

       5075 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2279] = !heapMem[localMem[2260]*6 + 6];
              ip = 5076;
      end

       5076 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2279] != 0 ? 5105 : 5077;
      end

       5077 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2280] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2280] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2280]] = 0;
              ip = 5078;
      end

       5078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 6] = localMem[2280];
              updateArrayLength(1, localMem[2276], 6);
              ip = 5079;
      end

       5079 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2281] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5080;
      end

       5080 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2282] = heapMem[localMem[2276]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5081;
      end

       5081 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2282] + 0 + i] = heapMem[NArea * localMem[2281] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2282], 0 + i);
                end
              end
              ip = 5082;
      end

       5082 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2283] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5083;
      end

       5083 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2284] = heapMem[localMem[2276]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5084;
      end

       5084 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2284] + 0 + i] = heapMem[NArea * localMem[2283] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2284], 0 + i);
                end
              end
              ip = 5085;
      end

       5085 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2285] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5086;
      end

       5086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2286] = heapMem[localMem[2276]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5087;
      end

       5087 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2287] = localMem[2273] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5088;
      end

       5088 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2287]) begin
                  heapMem[NArea * localMem[2286] + 0 + i] = heapMem[NArea * localMem[2285] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2286], 0 + i);
                end
              end
              ip = 5089;
      end

       5089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2288] = heapMem[localMem[2276]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5090;
      end

       5090 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2289] = localMem[2288] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5091;
      end

       5091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2290] = heapMem[localMem[2276]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5092;
      end

       5092 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5093;
      end

       5093 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2291] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5094;
      end

       5094 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5095;
      end

       5095 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2291] >= localMem[2289] ? 5101 : 5096;
      end

       5096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2292] = heapMem[localMem[2290]*6 + localMem[2291]];
              updateArrayLength(2, 0, 0);
              ip = 5097;
      end

       5097 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2292]*6 + 2] = localMem[2276];
              updateArrayLength(1, localMem[2292], 2);
              ip = 5098;
      end

       5098 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5099;
      end

       5099 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2291] = localMem[2291] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5100;
      end

       5100 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5094;
      end

       5101 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5102;
      end

       5102 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2293] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5103;
      end

       5103 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2293]] = localMem[2274];
              ip = 5104;
      end

       5104 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5112;
      end

       5105 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5106;
      end

       5106 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2294] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5107;
      end

       5107 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2295] = heapMem[localMem[2276]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5108;
      end

       5108 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2295] + 0 + i] = heapMem[NArea * localMem[2294] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2295], 0 + i);
                end
              end
              ip = 5109;
      end

       5109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2296] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5110;
      end

       5110 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2297] = heapMem[localMem[2276]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5111;
      end

       5111 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2297] + 0 + i] = heapMem[NArea * localMem[2296] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2297], 0 + i);
                end
              end
              ip = 5112;
      end

       5112 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5113;
      end

       5113 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2260]*6 + 0] = localMem[2273];
              updateArrayLength(1, localMem[2260], 0);
              ip = 5114;
      end

       5114 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*6 + 2] = localMem[2275];
              updateArrayLength(1, localMem[2276], 2);
              ip = 5115;
      end

       5115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2298] = heapMem[localMem[2275]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5116;
      end

       5116 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2299] = heapMem[localMem[2275]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5117;
      end

       5117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2300] = heapMem[localMem[2299]*6 + localMem[2298]];
              updateArrayLength(2, 0, 0);
              ip = 5118;
      end

       5118 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2300] != localMem[2260] ? 5137 : 5119;
      end

       5119 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2301] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5120;
      end

       5120 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2302] = heapMem[localMem[2301]*6 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5121;
      end

       5121 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2303] = heapMem[localMem[2275]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5122;
      end

       5122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2303]*6 + localMem[2298]] = localMem[2302];
              updateArrayLength(1, localMem[2303], localMem[2298]);
              ip = 5123;
      end

       5123 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2304] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5124;
      end

       5124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2305] = heapMem[localMem[2304]*6 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5125;
      end

       5125 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2306] = heapMem[localMem[2275]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5126;
      end

       5126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2306]*6 + localMem[2298]] = localMem[2305];
              updateArrayLength(1, localMem[2306], localMem[2298]);
              ip = 5127;
      end

       5127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2307] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5128;
      end

       5128 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2307]] = localMem[2273];
              ip = 5129;
      end

       5129 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2308] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5130;
      end

       5130 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2308]] = localMem[2273];
              ip = 5131;
      end

       5131 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2309] = localMem[2298] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5132;
      end

       5132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2275]*6 + 0] = localMem[2309];
              updateArrayLength(1, localMem[2275], 0);
              ip = 5133;
      end

       5133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2310] = heapMem[localMem[2275]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5134;
      end

       5134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2310]*6 + localMem[2309]] = localMem[2276];
              updateArrayLength(1, localMem[2310], localMem[2309]);
              ip = 5135;
      end

       5135 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5275;
      end

       5136 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5159;
      end

       5137 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5138;
      end

       5138 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 5139;
      end

       5139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2311] = heapMem[localMem[2275]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5140;
      end

       5140 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2312] = 0; k = arraySizes[localMem[2311]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2311] * NArea + i] == localMem[2260]) localMem[2312] = i + 1;
              end
              ip = 5141;
      end

       5141 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2312] = localMem[2312] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5142;
      end

       5142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2313] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5143;
      end

       5143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2314] = heapMem[localMem[2313]*6 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5144;
      end

       5144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2315] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5145;
      end

       5145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2316] = heapMem[localMem[2315]*6 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5146;
      end

       5146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2317] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5147;
      end

       5147 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2317]] = localMem[2273];
              ip = 5148;
      end

       5148 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2318] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5149;
      end

       5149 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2318]] = localMem[2273];
              ip = 5150;
      end

       5150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2319] = heapMem[localMem[2275]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5151;
      end

       5151 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2319] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2312], localMem[2319], arraySizes[localMem[2319]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2312] && i <= arraySizes[localMem[2319]]) begin
                  heapMem[NArea * localMem[2319] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2319] + localMem[2312]] = localMem[2314];                                    // Insert new value
              arraySizes[localMem[2319]] = arraySizes[localMem[2319]] + 1;                              // Increase array size
              ip = 5152;
      end

       5152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2320] = heapMem[localMem[2275]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5153;
      end

       5153 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2320] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2312], localMem[2320], arraySizes[localMem[2320]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2312] && i <= arraySizes[localMem[2320]]) begin
                  heapMem[NArea * localMem[2320] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2320] + localMem[2312]] = localMem[2316];                                    // Insert new value
              arraySizes[localMem[2320]] = arraySizes[localMem[2320]] + 1;                              // Increase array size
              ip = 5154;
      end

       5154 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2321] = heapMem[localMem[2275]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5155;
      end

       5155 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2322] = localMem[2312] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5156;
      end

       5156 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2321] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2322], localMem[2321], arraySizes[localMem[2321]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2322] && i <= arraySizes[localMem[2321]]) begin
                  heapMem[NArea * localMem[2321] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2321] + localMem[2322]] = localMem[2276];                                    // Insert new value
              arraySizes[localMem[2321]] = arraySizes[localMem[2321]] + 1;                              // Increase array size
              ip = 5157;
      end

       5157 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2275]*6 + 0] = heapMem[localMem[2275]*6 + 0] + 1;
              updateArrayLength(1, localMem[2275], 0);
              ip = 5158;
      end

       5158 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5275;
      end

       5159 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5160;
      end

       5160 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5161;
      end

       5161 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2323] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2323] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2323]] = 0;
              ip = 5162;
      end

       5162 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 0] = localMem[2273];
              updateArrayLength(1, localMem[2323], 0);
              ip = 5163;
      end

       5163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 2] = 0;
              updateArrayLength(1, localMem[2323], 2);
              ip = 5164;
      end

       5164 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2324] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2324] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2324]] = 0;
              ip = 5165;
      end

       5165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 4] = localMem[2324];
              updateArrayLength(1, localMem[2323], 4);
              ip = 5166;
      end

       5166 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2325] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2325] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2325]] = 0;
              ip = 5167;
      end

       5167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 5] = localMem[2325];
              updateArrayLength(1, localMem[2323], 5);
              ip = 5168;
      end

       5168 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 6] = 0;
              updateArrayLength(1, localMem[2323], 6);
              ip = 5169;
      end

       5169 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 3] = localMem[2271];
              updateArrayLength(1, localMem[2323], 3);
              ip = 5170;
      end

       5170 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2271]*6 + 1] = heapMem[localMem[2271]*6 + 1] + 1;
              updateArrayLength(1, localMem[2271], 1);
              ip = 5171;
      end

       5171 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 1] = heapMem[localMem[2271]*6 + 1];
              updateArrayLength(1, localMem[2323], 1);
              ip = 5172;
      end

       5172 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2326] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2326] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2326]] = 0;
              ip = 5173;
      end

       5173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 0] = localMem[2273];
              updateArrayLength(1, localMem[2326], 0);
              ip = 5174;
      end

       5174 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 2] = 0;
              updateArrayLength(1, localMem[2326], 2);
              ip = 5175;
      end

       5175 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2327] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2327] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2327]] = 0;
              ip = 5176;
      end

       5176 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 4] = localMem[2327];
              updateArrayLength(1, localMem[2326], 4);
              ip = 5177;
      end

       5177 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2328] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2328] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2328]] = 0;
              ip = 5178;
      end

       5178 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 5] = localMem[2328];
              updateArrayLength(1, localMem[2326], 5);
              ip = 5179;
      end

       5179 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 6] = 0;
              updateArrayLength(1, localMem[2326], 6);
              ip = 5180;
      end

       5180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 3] = localMem[2271];
              updateArrayLength(1, localMem[2326], 3);
              ip = 5181;
      end

       5181 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2271]*6 + 1] = heapMem[localMem[2271]*6 + 1] + 1;
              updateArrayLength(1, localMem[2271], 1);
              ip = 5182;
      end

       5182 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 1] = heapMem[localMem[2271]*6 + 1];
              updateArrayLength(1, localMem[2326], 1);
              ip = 5183;
      end

       5183 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2329] = !heapMem[localMem[2260]*6 + 6];
              ip = 5184;
      end

       5184 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2329] != 0 ? 5236 : 5185;
      end

       5185 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2330] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2330] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2330]] = 0;
              ip = 5186;
      end

       5186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 6] = localMem[2330];
              updateArrayLength(1, localMem[2323], 6);
              ip = 5187;
      end

       5187 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2331] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2331] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2331]] = 0;
              ip = 5188;
      end

       5188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 6] = localMem[2331];
              updateArrayLength(1, localMem[2326], 6);
              ip = 5189;
      end

       5189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2332] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5190;
      end

       5190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2333] = heapMem[localMem[2323]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5191;
      end

       5191 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2333] + 0 + i] = heapMem[NArea * localMem[2332] + 0 + i];
                  updateArrayLength(1, localMem[2333], 0 + i);
                end
              end
              ip = 5192;
      end

       5192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2334] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5193;
      end

       5193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2335] = heapMem[localMem[2323]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5194;
      end

       5194 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2335] + 0 + i] = heapMem[NArea * localMem[2334] + 0 + i];
                  updateArrayLength(1, localMem[2335], 0 + i);
                end
              end
              ip = 5195;
      end

       5195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2336] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5196;
      end

       5196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2337] = heapMem[localMem[2323]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5197;
      end

       5197 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2338] = localMem[2273] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5198;
      end

       5198 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2338]) begin
                  heapMem[NArea * localMem[2337] + 0 + i] = heapMem[NArea * localMem[2336] + 0 + i];
                  updateArrayLength(1, localMem[2337], 0 + i);
                end
              end
              ip = 5199;
      end

       5199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2339] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5200;
      end

       5200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2340] = heapMem[localMem[2326]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5201;
      end

       5201 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2340] + 0 + i] = heapMem[NArea * localMem[2339] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2340], 0 + i);
                end
              end
              ip = 5202;
      end

       5202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2341] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5203;
      end

       5203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2342] = heapMem[localMem[2326]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5204;
      end

       5204 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2342] + 0 + i] = heapMem[NArea * localMem[2341] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2342], 0 + i);
                end
              end
              ip = 5205;
      end

       5205 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2343] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5206;
      end

       5206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2344] = heapMem[localMem[2326]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5207;
      end

       5207 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2345] = localMem[2273] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5208;
      end

       5208 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2345]) begin
                  heapMem[NArea * localMem[2344] + 0 + i] = heapMem[NArea * localMem[2343] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2344], 0 + i);
                end
              end
              ip = 5209;
      end

       5209 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2346] = heapMem[localMem[2323]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5210;
      end

       5210 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2347] = localMem[2346] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5211;
      end

       5211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2348] = heapMem[localMem[2323]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5212;
      end

       5212 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5213;
      end

       5213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2349] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5214;
      end

       5214 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5215;
      end

       5215 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2349] >= localMem[2347] ? 5221 : 5216;
      end

       5216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2350] = heapMem[localMem[2348]*6 + localMem[2349]];
              updateArrayLength(2, 0, 0);
              ip = 5217;
      end

       5217 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2350]*6 + 2] = localMem[2323];
              updateArrayLength(1, localMem[2350], 2);
              ip = 5218;
      end

       5218 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5219;
      end

       5219 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2349] = localMem[2349] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5220;
      end

       5220 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5214;
      end

       5221 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5222;
      end

       5222 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2351] = heapMem[localMem[2326]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5223;
      end

       5223 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2352] = localMem[2351] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5224;
      end

       5224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2353] = heapMem[localMem[2326]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5225;
      end

       5225 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5226;
      end

       5226 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2354] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5227;
      end

       5227 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5228;
      end

       5228 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2354] >= localMem[2352] ? 5234 : 5229;
      end

       5229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2355] = heapMem[localMem[2353]*6 + localMem[2354]];
              updateArrayLength(2, 0, 0);
              ip = 5230;
      end

       5230 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2355]*6 + 2] = localMem[2326];
              updateArrayLength(1, localMem[2355], 2);
              ip = 5231;
      end

       5231 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5232;
      end

       5232 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2354] = localMem[2354] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5233;
      end

       5233 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5227;
      end

       5234 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5235;
      end

       5235 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5251;
      end

       5236 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5237;
      end

       5237 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2356] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2356] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2356]] = 0;
              ip = 5238;
      end

       5238 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2260]*6 + 6] = localMem[2356];
              updateArrayLength(1, localMem[2260], 6);
              ip = 5239;
      end

       5239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2357] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5240;
      end

       5240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2358] = heapMem[localMem[2323]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5241;
      end

       5241 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2358] + 0 + i] = heapMem[NArea * localMem[2357] + 0 + i];
                  updateArrayLength(1, localMem[2358], 0 + i);
                end
              end
              ip = 5242;
      end

       5242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2359] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5243;
      end

       5243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2360] = heapMem[localMem[2323]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5244;
      end

       5244 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2360] + 0 + i] = heapMem[NArea * localMem[2359] + 0 + i];
                  updateArrayLength(1, localMem[2360], 0 + i);
                end
              end
              ip = 5245;
      end

       5245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2361] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5246;
      end

       5246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2362] = heapMem[localMem[2326]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5247;
      end

       5247 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2362] + 0 + i] = heapMem[NArea * localMem[2361] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2362], 0 + i);
                end
              end
              ip = 5248;
      end

       5248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2363] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5249;
      end

       5249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2364] = heapMem[localMem[2326]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5250;
      end

       5250 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2364] + 0 + i] = heapMem[NArea * localMem[2363] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2364], 0 + i);
                end
              end
              ip = 5251;
      end

       5251 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5252;
      end

       5252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2323]*6 + 2] = localMem[2260];
              updateArrayLength(1, localMem[2323], 2);
              ip = 5253;
      end

       5253 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2326]*6 + 2] = localMem[2260];
              updateArrayLength(1, localMem[2326], 2);
              ip = 5254;
      end

       5254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2365] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5255;
      end

       5255 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2366] = heapMem[localMem[2365]*6 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5256;
      end

       5256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2367] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5257;
      end

       5257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2368] = heapMem[localMem[2367]*6 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5258;
      end

       5258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2369] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5259;
      end

       5259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2369]*6 + 0] = localMem[2366];
              updateArrayLength(1, localMem[2369], 0);
              ip = 5260;
      end

       5260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2370] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5261;
      end

       5261 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2370]*6 + 0] = localMem[2368];
              updateArrayLength(1, localMem[2370], 0);
              ip = 5262;
      end

       5262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2371] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5263;
      end

       5263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2371]*6 + 0] = localMem[2323];
              updateArrayLength(1, localMem[2371], 0);
              ip = 5264;
      end

       5264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2372] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5265;
      end

       5265 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2372]*6 + 1] = localMem[2326];
              updateArrayLength(1, localMem[2372], 1);
              ip = 5266;
      end

       5266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2260]*6 + 0] = 1;
              updateArrayLength(1, localMem[2260], 0);
              ip = 5267;
      end

       5267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2373] = heapMem[localMem[2260]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5268;
      end

       5268 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2373]] = 1;
              ip = 5269;
      end

       5269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2374] = heapMem[localMem[2260]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5270;
      end

       5270 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2374]] = 1;
              ip = 5271;
      end

       5271 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2375] = heapMem[localMem[2260]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5272;
      end

       5272 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2375]] = 2;
              ip = 5273;
      end

       5273 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5275;
      end

       5274 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5280;
      end

       5275 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5276;
      end

       5276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2269] = 1;
              updateArrayLength(2, 0, 0);
              ip = 5277;
      end

       5277 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5280;
      end

       5278 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5279;
      end

       5279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2269] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5280;
      end

       5280 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5281;
      end

       5281 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5282;
      end

       5282 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5283;
      end

       5283 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5284;
      end

       5284 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[1901]] = 0;
              freedArrays[freedArraysTop] = localMem[1901];
              freedArraysTop = freedArraysTop + 1;
              ip = 5285;
      end

       5285 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2376] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2376] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2376]] = 0;
              ip = 5286;
      end

       5286 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5287;
      end

       5287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2377] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5288;
      end

       5288 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2377] != 0 ? 5311 : 5289;
      end

       5289 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2378] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2378] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2378]] = 0;
              ip = 5290;
      end

       5290 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 0] = 1;
              updateArrayLength(1, localMem[2378], 0);
              ip = 5291;
      end

       5291 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 2] = 0;
              updateArrayLength(1, localMem[2378], 2);
              ip = 5292;
      end

       5292 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2379] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2379] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2379]] = 0;
              ip = 5293;
      end

       5293 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 4] = localMem[2379];
              updateArrayLength(1, localMem[2378], 4);
              ip = 5294;
      end

       5294 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2380] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2380] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2380]] = 0;
              ip = 5295;
      end

       5295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 5] = localMem[2380];
              updateArrayLength(1, localMem[2378], 5);
              ip = 5296;
      end

       5296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 6] = 0;
              updateArrayLength(1, localMem[2378], 6);
              ip = 5297;
      end

       5297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 3] = localMem[0];
              updateArrayLength(1, localMem[2378], 3);
              ip = 5298;
      end

       5298 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 1] = heapMem[localMem[0]*6 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 5299;
      end

       5299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2378]*6 + 1] = heapMem[localMem[0]*6 + 1];
              updateArrayLength(1, localMem[2378], 1);
              ip = 5300;
      end

       5300 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2381] = heapMem[localMem[2378]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5301;
      end

       5301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2381]*6 + 0] = 6;
              updateArrayLength(1, localMem[2381], 0);
              ip = 5302;
      end

       5302 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2382] = heapMem[localMem[2378]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5303;
      end

       5303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2382]*6 + 0] = 66;
              updateArrayLength(1, localMem[2382], 0);
              ip = 5304;
      end

       5304 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 5305;
      end

       5305 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*6 + 3] = localMem[2378];
              updateArrayLength(1, localMem[0], 3);
              ip = 5306;
      end

       5306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2383] = heapMem[localMem[2378]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5307;
      end

       5307 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2383]] = 1;
              ip = 5308;
      end

       5308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2384] = heapMem[localMem[2378]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5309;
      end

       5309 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2384]] = 1;
              ip = 5310;
      end

       5310 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6339;
      end

       5311 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5312;
      end

       5312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2385] = heapMem[localMem[2377]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5313;
      end

       5313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2386] = heapMem[localMem[0]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5314;
      end

       5314 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2385] >= localMem[2386] ? 5350 : 5315;
      end

       5315 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2387] = heapMem[localMem[2377]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5316;
      end

       5316 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2387] != 0 ? 5349 : 5317;
      end

       5317 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2388] = !heapMem[localMem[2377]*6 + 6];
              ip = 5318;
      end

       5318 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2388] == 0 ? 5348 : 5319;
      end

       5319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2389] = heapMem[localMem[2377]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5320;
      end

       5320 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2390] = 0; k = arraySizes[localMem[2389]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2389] * NArea + i] == 6) localMem[2390] = i + 1;
              end
              ip = 5321;
      end

       5321 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2390] == 0 ? 5326 : 5322;
      end

       5322 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2390] = localMem[2390] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5323;
      end

       5323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2391] = heapMem[localMem[2377]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5324;
      end

       5324 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2391]*6 + localMem[2390]] = 66;
              updateArrayLength(1, localMem[2391], localMem[2390]);
              ip = 5325;
      end

       5325 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6339;
      end

       5326 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5327;
      end

       5327 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2389]] = localMem[2385];
              ip = 5328;
      end

       5328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2392] = heapMem[localMem[2377]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5329;
      end

       5329 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2392]] = localMem[2385];
              ip = 5330;
      end

       5330 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[2389]];
//$display("AAAAA k=%d  source2=%d", k, 6);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[2389] * NArea + i]);
                if (i < k && heapMem[localMem[2389] * NArea + i] > 6) j = j + 1;
              end
              localMem[2393] = j;
              ip = 5331;
      end

       5331 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2393] != 0 ? 5339 : 5332;
      end

       5332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2394] = heapMem[localMem[2377]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5333;
      end

       5333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2394]*6 + localMem[2385]] = 6;
              updateArrayLength(1, localMem[2394], localMem[2385]);
              ip = 5334;
      end

       5334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2395] = heapMem[localMem[2377]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5335;
      end

       5335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2395]*6 + localMem[2385]] = 66;
              updateArrayLength(1, localMem[2395], localMem[2385]);
              ip = 5336;
      end

       5336 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2377]*6 + 0] = localMem[2385] + 1;
              updateArrayLength(1, localMem[2377], 0);
              ip = 5337;
      end

       5337 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 5338;
      end

       5338 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6339;
      end

       5339 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5340;
      end

       5340 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[2389]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2389] * NArea + i] < 6) j = j + 1;
              end
              localMem[2396] = j;
              ip = 5341;
      end

       5341 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2397] = heapMem[localMem[2377]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5342;
      end

       5342 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2397] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2396], localMem[2397], arraySizes[localMem[2397]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2396] && i <= arraySizes[localMem[2397]]) begin
                  heapMem[NArea * localMem[2397] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2397] + localMem[2396]] = 6;                                    // Insert new value
              arraySizes[localMem[2397]] = arraySizes[localMem[2397]] + 1;                              // Increase array size
              ip = 5343;
      end

       5343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2398] = heapMem[localMem[2377]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5344;
      end

       5344 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2398] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2396], localMem[2398], arraySizes[localMem[2398]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2396] && i <= arraySizes[localMem[2398]]) begin
                  heapMem[NArea * localMem[2398] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2398] + localMem[2396]] = 66;                                    // Insert new value
              arraySizes[localMem[2398]] = arraySizes[localMem[2398]] + 1;                              // Increase array size
              ip = 5345;
      end

       5345 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2377]*6 + 0] = heapMem[localMem[2377]*6 + 0] + 1;
              updateArrayLength(1, localMem[2377], 0);
              ip = 5346;
      end

       5346 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 5347;
      end

       5347 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6339;
      end

       5348 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5349;
      end

       5349 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5350;
      end

       5350 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5351;
      end

       5351 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2399] = heapMem[localMem[0]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5352;
      end

       5352 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5353;
      end

       5353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2401] = heapMem[localMem[2399]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5354;
      end

       5354 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2402] = heapMem[localMem[2399]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5355;
      end

       5355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2403] = heapMem[localMem[2402]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5356;
      end

       5356 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2401] <  localMem[2403] ? 5576 : 5357;
      end

       5357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2404] = localMem[2403];
              updateArrayLength(2, 0, 0);
              ip = 5358;
      end

       5358 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2404] = localMem[2404] >> 1;
              ip = 5359;
      end

       5359 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2405] = localMem[2404] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5360;
      end

       5360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2406] = heapMem[localMem[2399]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5361;
      end

       5361 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2406] == 0 ? 5458 : 5362;
      end

       5362 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2407] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2407] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2407]] = 0;
              ip = 5363;
      end

       5363 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 0] = localMem[2404];
              updateArrayLength(1, localMem[2407], 0);
              ip = 5364;
      end

       5364 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 2] = 0;
              updateArrayLength(1, localMem[2407], 2);
              ip = 5365;
      end

       5365 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2408] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2408] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2408]] = 0;
              ip = 5366;
      end

       5366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 4] = localMem[2408];
              updateArrayLength(1, localMem[2407], 4);
              ip = 5367;
      end

       5367 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2409] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2409] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2409]] = 0;
              ip = 5368;
      end

       5368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 5] = localMem[2409];
              updateArrayLength(1, localMem[2407], 5);
              ip = 5369;
      end

       5369 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 6] = 0;
              updateArrayLength(1, localMem[2407], 6);
              ip = 5370;
      end

       5370 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 3] = localMem[2402];
              updateArrayLength(1, localMem[2407], 3);
              ip = 5371;
      end

       5371 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2402]*6 + 1] = heapMem[localMem[2402]*6 + 1] + 1;
              updateArrayLength(1, localMem[2402], 1);
              ip = 5372;
      end

       5372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 1] = heapMem[localMem[2402]*6 + 1];
              updateArrayLength(1, localMem[2407], 1);
              ip = 5373;
      end

       5373 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2410] = !heapMem[localMem[2399]*6 + 6];
              ip = 5374;
      end

       5374 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2410] != 0 ? 5403 : 5375;
      end

       5375 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2411] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2411] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2411]] = 0;
              ip = 5376;
      end

       5376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 6] = localMem[2411];
              updateArrayLength(1, localMem[2407], 6);
              ip = 5377;
      end

       5377 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2412] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5378;
      end

       5378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2413] = heapMem[localMem[2407]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5379;
      end

       5379 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2413] + 0 + i] = heapMem[NArea * localMem[2412] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2413], 0 + i);
                end
              end
              ip = 5380;
      end

       5380 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2414] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5381;
      end

       5381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2415] = heapMem[localMem[2407]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5382;
      end

       5382 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2415] + 0 + i] = heapMem[NArea * localMem[2414] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2415], 0 + i);
                end
              end
              ip = 5383;
      end

       5383 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2416] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5384;
      end

       5384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2417] = heapMem[localMem[2407]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5385;
      end

       5385 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2418] = localMem[2404] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5386;
      end

       5386 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2418]) begin
                  heapMem[NArea * localMem[2417] + 0 + i] = heapMem[NArea * localMem[2416] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2417], 0 + i);
                end
              end
              ip = 5387;
      end

       5387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2419] = heapMem[localMem[2407]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5388;
      end

       5388 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2420] = localMem[2419] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5389;
      end

       5389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2421] = heapMem[localMem[2407]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5390;
      end

       5390 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5391;
      end

       5391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2422] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5392;
      end

       5392 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5393;
      end

       5393 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2422] >= localMem[2420] ? 5399 : 5394;
      end

       5394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2423] = heapMem[localMem[2421]*6 + localMem[2422]];
              updateArrayLength(2, 0, 0);
              ip = 5395;
      end

       5395 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2423]*6 + 2] = localMem[2407];
              updateArrayLength(1, localMem[2423], 2);
              ip = 5396;
      end

       5396 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5397;
      end

       5397 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2422] = localMem[2422] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5398;
      end

       5398 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5392;
      end

       5399 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5400;
      end

       5400 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2424] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5401;
      end

       5401 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2424]] = localMem[2405];
              ip = 5402;
      end

       5402 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5410;
      end

       5403 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5404;
      end

       5404 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2425] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5405;
      end

       5405 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2426] = heapMem[localMem[2407]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5406;
      end

       5406 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2426] + 0 + i] = heapMem[NArea * localMem[2425] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2426], 0 + i);
                end
              end
              ip = 5407;
      end

       5407 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2427] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5408;
      end

       5408 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2428] = heapMem[localMem[2407]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5409;
      end

       5409 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2428] + 0 + i] = heapMem[NArea * localMem[2427] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2428], 0 + i);
                end
              end
              ip = 5410;
      end

       5410 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5411;
      end

       5411 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2399]*6 + 0] = localMem[2404];
              updateArrayLength(1, localMem[2399], 0);
              ip = 5412;
      end

       5412 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2407]*6 + 2] = localMem[2406];
              updateArrayLength(1, localMem[2407], 2);
              ip = 5413;
      end

       5413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2429] = heapMem[localMem[2406]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5414;
      end

       5414 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2430] = heapMem[localMem[2406]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5415;
      end

       5415 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2431] = heapMem[localMem[2430]*6 + localMem[2429]];
              updateArrayLength(2, 0, 0);
              ip = 5416;
      end

       5416 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2431] != localMem[2399] ? 5435 : 5417;
      end

       5417 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2432] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5418;
      end

       5418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2433] = heapMem[localMem[2432]*6 + localMem[2404]];
              updateArrayLength(2, 0, 0);
              ip = 5419;
      end

       5419 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2434] = heapMem[localMem[2406]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5420;
      end

       5420 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2434]*6 + localMem[2429]] = localMem[2433];
              updateArrayLength(1, localMem[2434], localMem[2429]);
              ip = 5421;
      end

       5421 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2435] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5422;
      end

       5422 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2436] = heapMem[localMem[2435]*6 + localMem[2404]];
              updateArrayLength(2, 0, 0);
              ip = 5423;
      end

       5423 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2437] = heapMem[localMem[2406]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5424;
      end

       5424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2437]*6 + localMem[2429]] = localMem[2436];
              updateArrayLength(1, localMem[2437], localMem[2429]);
              ip = 5425;
      end

       5425 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2438] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5426;
      end

       5426 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2438]] = localMem[2404];
              ip = 5427;
      end

       5427 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2439] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5428;
      end

       5428 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2439]] = localMem[2404];
              ip = 5429;
      end

       5429 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2440] = localMem[2429] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5430;
      end

       5430 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2406]*6 + 0] = localMem[2440];
              updateArrayLength(1, localMem[2406], 0);
              ip = 5431;
      end

       5431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2441] = heapMem[localMem[2406]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5432;
      end

       5432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2441]*6 + localMem[2440]] = localMem[2407];
              updateArrayLength(1, localMem[2441], localMem[2440]);
              ip = 5433;
      end

       5433 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5573;
      end

       5434 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5457;
      end

       5435 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5436;
      end

       5436 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 5437;
      end

       5437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2442] = heapMem[localMem[2406]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5438;
      end

       5438 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2443] = 0; k = arraySizes[localMem[2442]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2442] * NArea + i] == localMem[2399]) localMem[2443] = i + 1;
              end
              ip = 5439;
      end

       5439 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2443] = localMem[2443] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5440;
      end

       5440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2444] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5441;
      end

       5441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2445] = heapMem[localMem[2444]*6 + localMem[2404]];
              updateArrayLength(2, 0, 0);
              ip = 5442;
      end

       5442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2446] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5443;
      end

       5443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2447] = heapMem[localMem[2446]*6 + localMem[2404]];
              updateArrayLength(2, 0, 0);
              ip = 5444;
      end

       5444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2448] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5445;
      end

       5445 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2448]] = localMem[2404];
              ip = 5446;
      end

       5446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2449] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5447;
      end

       5447 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2449]] = localMem[2404];
              ip = 5448;
      end

       5448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2450] = heapMem[localMem[2406]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5449;
      end

       5449 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2450] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2443], localMem[2450], arraySizes[localMem[2450]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2443] && i <= arraySizes[localMem[2450]]) begin
                  heapMem[NArea * localMem[2450] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2450] + localMem[2443]] = localMem[2445];                                    // Insert new value
              arraySizes[localMem[2450]] = arraySizes[localMem[2450]] + 1;                              // Increase array size
              ip = 5450;
      end

       5450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2451] = heapMem[localMem[2406]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5451;
      end

       5451 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2451] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2443], localMem[2451], arraySizes[localMem[2451]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2443] && i <= arraySizes[localMem[2451]]) begin
                  heapMem[NArea * localMem[2451] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2451] + localMem[2443]] = localMem[2447];                                    // Insert new value
              arraySizes[localMem[2451]] = arraySizes[localMem[2451]] + 1;                              // Increase array size
              ip = 5452;
      end

       5452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2452] = heapMem[localMem[2406]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5453;
      end

       5453 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2453] = localMem[2443] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5454;
      end

       5454 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2452] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2453], localMem[2452], arraySizes[localMem[2452]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2453] && i <= arraySizes[localMem[2452]]) begin
                  heapMem[NArea * localMem[2452] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2452] + localMem[2453]] = localMem[2407];                                    // Insert new value
              arraySizes[localMem[2452]] = arraySizes[localMem[2452]] + 1;                              // Increase array size
              ip = 5455;
      end

       5455 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2406]*6 + 0] = heapMem[localMem[2406]*6 + 0] + 1;
              updateArrayLength(1, localMem[2406], 0);
              ip = 5456;
      end

       5456 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5573;
      end

       5457 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5458;
      end

       5458 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5459;
      end

       5459 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2454] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2454] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2454]] = 0;
              ip = 5460;
      end

       5460 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 0] = localMem[2404];
              updateArrayLength(1, localMem[2454], 0);
              ip = 5461;
      end

       5461 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 2] = 0;
              updateArrayLength(1, localMem[2454], 2);
              ip = 5462;
      end

       5462 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2455] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2455] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2455]] = 0;
              ip = 5463;
      end

       5463 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 4] = localMem[2455];
              updateArrayLength(1, localMem[2454], 4);
              ip = 5464;
      end

       5464 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2456] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2456] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2456]] = 0;
              ip = 5465;
      end

       5465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 5] = localMem[2456];
              updateArrayLength(1, localMem[2454], 5);
              ip = 5466;
      end

       5466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 6] = 0;
              updateArrayLength(1, localMem[2454], 6);
              ip = 5467;
      end

       5467 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 3] = localMem[2402];
              updateArrayLength(1, localMem[2454], 3);
              ip = 5468;
      end

       5468 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2402]*6 + 1] = heapMem[localMem[2402]*6 + 1] + 1;
              updateArrayLength(1, localMem[2402], 1);
              ip = 5469;
      end

       5469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 1] = heapMem[localMem[2402]*6 + 1];
              updateArrayLength(1, localMem[2454], 1);
              ip = 5470;
      end

       5470 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2457] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2457] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2457]] = 0;
              ip = 5471;
      end

       5471 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 0] = localMem[2404];
              updateArrayLength(1, localMem[2457], 0);
              ip = 5472;
      end

       5472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 2] = 0;
              updateArrayLength(1, localMem[2457], 2);
              ip = 5473;
      end

       5473 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2458] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2458] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2458]] = 0;
              ip = 5474;
      end

       5474 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 4] = localMem[2458];
              updateArrayLength(1, localMem[2457], 4);
              ip = 5475;
      end

       5475 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2459] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2459] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2459]] = 0;
              ip = 5476;
      end

       5476 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 5] = localMem[2459];
              updateArrayLength(1, localMem[2457], 5);
              ip = 5477;
      end

       5477 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 6] = 0;
              updateArrayLength(1, localMem[2457], 6);
              ip = 5478;
      end

       5478 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 3] = localMem[2402];
              updateArrayLength(1, localMem[2457], 3);
              ip = 5479;
      end

       5479 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2402]*6 + 1] = heapMem[localMem[2402]*6 + 1] + 1;
              updateArrayLength(1, localMem[2402], 1);
              ip = 5480;
      end

       5480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 1] = heapMem[localMem[2402]*6 + 1];
              updateArrayLength(1, localMem[2457], 1);
              ip = 5481;
      end

       5481 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2460] = !heapMem[localMem[2399]*6 + 6];
              ip = 5482;
      end

       5482 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2460] != 0 ? 5534 : 5483;
      end

       5483 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2461] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2461] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2461]] = 0;
              ip = 5484;
      end

       5484 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 6] = localMem[2461];
              updateArrayLength(1, localMem[2454], 6);
              ip = 5485;
      end

       5485 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2462] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2462] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2462]] = 0;
              ip = 5486;
      end

       5486 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 6] = localMem[2462];
              updateArrayLength(1, localMem[2457], 6);
              ip = 5487;
      end

       5487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2463] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5488;
      end

       5488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2464] = heapMem[localMem[2454]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5489;
      end

       5489 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2464] + 0 + i] = heapMem[NArea * localMem[2463] + 0 + i];
                  updateArrayLength(1, localMem[2464], 0 + i);
                end
              end
              ip = 5490;
      end

       5490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2465] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5491;
      end

       5491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2466] = heapMem[localMem[2454]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5492;
      end

       5492 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2466] + 0 + i] = heapMem[NArea * localMem[2465] + 0 + i];
                  updateArrayLength(1, localMem[2466], 0 + i);
                end
              end
              ip = 5493;
      end

       5493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2467] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5494;
      end

       5494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2468] = heapMem[localMem[2454]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5495;
      end

       5495 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2469] = localMem[2404] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5496;
      end

       5496 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2469]) begin
                  heapMem[NArea * localMem[2468] + 0 + i] = heapMem[NArea * localMem[2467] + 0 + i];
                  updateArrayLength(1, localMem[2468], 0 + i);
                end
              end
              ip = 5497;
      end

       5497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2470] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5498;
      end

       5498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2471] = heapMem[localMem[2457]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5499;
      end

       5499 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2471] + 0 + i] = heapMem[NArea * localMem[2470] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2471], 0 + i);
                end
              end
              ip = 5500;
      end

       5500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2472] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5501;
      end

       5501 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2473] = heapMem[localMem[2457]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5502;
      end

       5502 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2473] + 0 + i] = heapMem[NArea * localMem[2472] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2473], 0 + i);
                end
              end
              ip = 5503;
      end

       5503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2474] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5504;
      end

       5504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2475] = heapMem[localMem[2457]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5505;
      end

       5505 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2476] = localMem[2404] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5506;
      end

       5506 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2476]) begin
                  heapMem[NArea * localMem[2475] + 0 + i] = heapMem[NArea * localMem[2474] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2475], 0 + i);
                end
              end
              ip = 5507;
      end

       5507 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2477] = heapMem[localMem[2454]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5508;
      end

       5508 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2478] = localMem[2477] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5509;
      end

       5509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2479] = heapMem[localMem[2454]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5510;
      end

       5510 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5511;
      end

       5511 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2480] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5512;
      end

       5512 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5513;
      end

       5513 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2480] >= localMem[2478] ? 5519 : 5514;
      end

       5514 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2481] = heapMem[localMem[2479]*6 + localMem[2480]];
              updateArrayLength(2, 0, 0);
              ip = 5515;
      end

       5515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2481]*6 + 2] = localMem[2454];
              updateArrayLength(1, localMem[2481], 2);
              ip = 5516;
      end

       5516 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5517;
      end

       5517 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2480] = localMem[2480] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5518;
      end

       5518 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5512;
      end

       5519 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5520;
      end

       5520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2482] = heapMem[localMem[2457]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5521;
      end

       5521 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2483] = localMem[2482] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5522;
      end

       5522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2484] = heapMem[localMem[2457]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5523;
      end

       5523 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5524;
      end

       5524 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2485] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5525;
      end

       5525 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5526;
      end

       5526 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2485] >= localMem[2483] ? 5532 : 5527;
      end

       5527 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2486] = heapMem[localMem[2484]*6 + localMem[2485]];
              updateArrayLength(2, 0, 0);
              ip = 5528;
      end

       5528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2486]*6 + 2] = localMem[2457];
              updateArrayLength(1, localMem[2486], 2);
              ip = 5529;
      end

       5529 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5530;
      end

       5530 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2485] = localMem[2485] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5531;
      end

       5531 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5525;
      end

       5532 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5533;
      end

       5533 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5549;
      end

       5534 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5535;
      end

       5535 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2487] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2487] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2487]] = 0;
              ip = 5536;
      end

       5536 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2399]*6 + 6] = localMem[2487];
              updateArrayLength(1, localMem[2399], 6);
              ip = 5537;
      end

       5537 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2488] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5538;
      end

       5538 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2489] = heapMem[localMem[2454]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5539;
      end

       5539 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2489] + 0 + i] = heapMem[NArea * localMem[2488] + 0 + i];
                  updateArrayLength(1, localMem[2489], 0 + i);
                end
              end
              ip = 5540;
      end

       5540 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2490] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5541;
      end

       5541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2491] = heapMem[localMem[2454]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5542;
      end

       5542 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2491] + 0 + i] = heapMem[NArea * localMem[2490] + 0 + i];
                  updateArrayLength(1, localMem[2491], 0 + i);
                end
              end
              ip = 5543;
      end

       5543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2492] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5544;
      end

       5544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2493] = heapMem[localMem[2457]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5545;
      end

       5545 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2493] + 0 + i] = heapMem[NArea * localMem[2492] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2493], 0 + i);
                end
              end
              ip = 5546;
      end

       5546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2494] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5547;
      end

       5547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2495] = heapMem[localMem[2457]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5548;
      end

       5548 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2404]) begin
                  heapMem[NArea * localMem[2495] + 0 + i] = heapMem[NArea * localMem[2494] + localMem[2405] + i];
                  updateArrayLength(1, localMem[2495], 0 + i);
                end
              end
              ip = 5549;
      end

       5549 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5550;
      end

       5550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2454]*6 + 2] = localMem[2399];
              updateArrayLength(1, localMem[2454], 2);
              ip = 5551;
      end

       5551 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2457]*6 + 2] = localMem[2399];
              updateArrayLength(1, localMem[2457], 2);
              ip = 5552;
      end

       5552 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2496] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5553;
      end

       5553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2497] = heapMem[localMem[2496]*6 + localMem[2404]];
              updateArrayLength(2, 0, 0);
              ip = 5554;
      end

       5554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2498] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5555;
      end

       5555 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2499] = heapMem[localMem[2498]*6 + localMem[2404]];
              updateArrayLength(2, 0, 0);
              ip = 5556;
      end

       5556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2500] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5557;
      end

       5557 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2500]*6 + 0] = localMem[2497];
              updateArrayLength(1, localMem[2500], 0);
              ip = 5558;
      end

       5558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2501] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5559;
      end

       5559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2501]*6 + 0] = localMem[2499];
              updateArrayLength(1, localMem[2501], 0);
              ip = 5560;
      end

       5560 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2502] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5561;
      end

       5561 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2502]*6 + 0] = localMem[2454];
              updateArrayLength(1, localMem[2502], 0);
              ip = 5562;
      end

       5562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2503] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5563;
      end

       5563 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2503]*6 + 1] = localMem[2457];
              updateArrayLength(1, localMem[2503], 1);
              ip = 5564;
      end

       5564 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2399]*6 + 0] = 1;
              updateArrayLength(1, localMem[2399], 0);
              ip = 5565;
      end

       5565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2504] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5566;
      end

       5566 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2504]] = 1;
              ip = 5567;
      end

       5567 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2505] = heapMem[localMem[2399]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5568;
      end

       5568 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2505]] = 1;
              ip = 5569;
      end

       5569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2506] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5570;
      end

       5570 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2506]] = 2;
              ip = 5571;
      end

       5571 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5573;
      end

       5572 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5578;
      end

       5573 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5574;
      end

       5574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2400] = 1;
              updateArrayLength(2, 0, 0);
              ip = 5575;
      end

       5575 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5578;
      end

       5576 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5577;
      end

       5577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2400] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5578;
      end

       5578 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5579;
      end

       5579 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5580;
      end

       5580 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5581;
      end

       5581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2507] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5582;
      end

       5582 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5583;
      end

       5583 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2507] >= 99 ? 6081 : 5584;
      end

       5584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2508] = heapMem[localMem[2399]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5585;
      end

       5585 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2509] = localMem[2508] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5586;
      end

       5586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2510] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5587;
      end

       5587 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2511] = heapMem[localMem[2510]*6 + localMem[2509]];
              updateArrayLength(2, 0, 0);
              ip = 5588;
      end

       5588 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 6 <= localMem[2511] ? 5829 : 5589;
      end

       5589 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2512] = !heapMem[localMem[2399]*6 + 6];
              ip = 5590;
      end

       5590 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2512] == 0 ? 5595 : 5591;
      end

       5591 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 0] = localMem[2399];
              updateArrayLength(1, localMem[2376], 0);
              ip = 5592;
      end

       5592 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 1] = 2;
              updateArrayLength(1, localMem[2376], 1);
              ip = 5593;
      end

       5593 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[2376]*6 + 2] = localMem[2508] - 1;
              updateArrayLength(1, localMem[2376], 2);
              ip = 5594;
      end

       5594 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6085;
      end

       5595 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5596;
      end

       5596 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2513] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5597;
      end

       5597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2514] = heapMem[localMem[2513]*6 + localMem[2508]];
              updateArrayLength(2, 0, 0);
              ip = 5598;
      end

       5598 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5599;
      end

       5599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2516] = heapMem[localMem[2514]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5600;
      end

       5600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2517] = heapMem[localMem[2514]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5601;
      end

       5601 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2518] = heapMem[localMem[2517]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5602;
      end

       5602 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2516] <  localMem[2518] ? 5822 : 5603;
      end

       5603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2519] = localMem[2518];
              updateArrayLength(2, 0, 0);
              ip = 5604;
      end

       5604 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2519] = localMem[2519] >> 1;
              ip = 5605;
      end

       5605 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2520] = localMem[2519] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5606;
      end

       5606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2521] = heapMem[localMem[2514]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5607;
      end

       5607 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2521] == 0 ? 5704 : 5608;
      end

       5608 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2522] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2522] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2522]] = 0;
              ip = 5609;
      end

       5609 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 0] = localMem[2519];
              updateArrayLength(1, localMem[2522], 0);
              ip = 5610;
      end

       5610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 2] = 0;
              updateArrayLength(1, localMem[2522], 2);
              ip = 5611;
      end

       5611 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2523] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2523] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2523]] = 0;
              ip = 5612;
      end

       5612 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 4] = localMem[2523];
              updateArrayLength(1, localMem[2522], 4);
              ip = 5613;
      end

       5613 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2524] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2524] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2524]] = 0;
              ip = 5614;
      end

       5614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 5] = localMem[2524];
              updateArrayLength(1, localMem[2522], 5);
              ip = 5615;
      end

       5615 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 6] = 0;
              updateArrayLength(1, localMem[2522], 6);
              ip = 5616;
      end

       5616 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 3] = localMem[2517];
              updateArrayLength(1, localMem[2522], 3);
              ip = 5617;
      end

       5617 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2517]*6 + 1] = heapMem[localMem[2517]*6 + 1] + 1;
              updateArrayLength(1, localMem[2517], 1);
              ip = 5618;
      end

       5618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 1] = heapMem[localMem[2517]*6 + 1];
              updateArrayLength(1, localMem[2522], 1);
              ip = 5619;
      end

       5619 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2525] = !heapMem[localMem[2514]*6 + 6];
              ip = 5620;
      end

       5620 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2525] != 0 ? 5649 : 5621;
      end

       5621 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2526] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2526] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2526]] = 0;
              ip = 5622;
      end

       5622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 6] = localMem[2526];
              updateArrayLength(1, localMem[2522], 6);
              ip = 5623;
      end

       5623 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2527] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5624;
      end

       5624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2528] = heapMem[localMem[2522]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5625;
      end

       5625 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2528] + 0 + i] = heapMem[NArea * localMem[2527] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2528], 0 + i);
                end
              end
              ip = 5626;
      end

       5626 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2529] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5627;
      end

       5627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2530] = heapMem[localMem[2522]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5628;
      end

       5628 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2530] + 0 + i] = heapMem[NArea * localMem[2529] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2530], 0 + i);
                end
              end
              ip = 5629;
      end

       5629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2531] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5630;
      end

       5630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2532] = heapMem[localMem[2522]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5631;
      end

       5631 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2533] = localMem[2519] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5632;
      end

       5632 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2533]) begin
                  heapMem[NArea * localMem[2532] + 0 + i] = heapMem[NArea * localMem[2531] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2532], 0 + i);
                end
              end
              ip = 5633;
      end

       5633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2534] = heapMem[localMem[2522]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5634;
      end

       5634 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2535] = localMem[2534] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5635;
      end

       5635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2536] = heapMem[localMem[2522]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5636;
      end

       5636 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5637;
      end

       5637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2537] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5638;
      end

       5638 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5639;
      end

       5639 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2537] >= localMem[2535] ? 5645 : 5640;
      end

       5640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2538] = heapMem[localMem[2536]*6 + localMem[2537]];
              updateArrayLength(2, 0, 0);
              ip = 5641;
      end

       5641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2538]*6 + 2] = localMem[2522];
              updateArrayLength(1, localMem[2538], 2);
              ip = 5642;
      end

       5642 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5643;
      end

       5643 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2537] = localMem[2537] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5644;
      end

       5644 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5638;
      end

       5645 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5646;
      end

       5646 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2539] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5647;
      end

       5647 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2539]] = localMem[2520];
              ip = 5648;
      end

       5648 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5656;
      end

       5649 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5650;
      end

       5650 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2540] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5651;
      end

       5651 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2541] = heapMem[localMem[2522]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5652;
      end

       5652 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2541] + 0 + i] = heapMem[NArea * localMem[2540] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2541], 0 + i);
                end
              end
              ip = 5653;
      end

       5653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2542] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5654;
      end

       5654 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2543] = heapMem[localMem[2522]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5655;
      end

       5655 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2543] + 0 + i] = heapMem[NArea * localMem[2542] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2543], 0 + i);
                end
              end
              ip = 5656;
      end

       5656 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5657;
      end

       5657 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2514]*6 + 0] = localMem[2519];
              updateArrayLength(1, localMem[2514], 0);
              ip = 5658;
      end

       5658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2522]*6 + 2] = localMem[2521];
              updateArrayLength(1, localMem[2522], 2);
              ip = 5659;
      end

       5659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2544] = heapMem[localMem[2521]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5660;
      end

       5660 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2545] = heapMem[localMem[2521]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5661;
      end

       5661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2546] = heapMem[localMem[2545]*6 + localMem[2544]];
              updateArrayLength(2, 0, 0);
              ip = 5662;
      end

       5662 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2546] != localMem[2514] ? 5681 : 5663;
      end

       5663 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2547] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5664;
      end

       5664 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2548] = heapMem[localMem[2547]*6 + localMem[2519]];
              updateArrayLength(2, 0, 0);
              ip = 5665;
      end

       5665 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2549] = heapMem[localMem[2521]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5666;
      end

       5666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2549]*6 + localMem[2544]] = localMem[2548];
              updateArrayLength(1, localMem[2549], localMem[2544]);
              ip = 5667;
      end

       5667 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2550] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5668;
      end

       5668 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2551] = heapMem[localMem[2550]*6 + localMem[2519]];
              updateArrayLength(2, 0, 0);
              ip = 5669;
      end

       5669 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2552] = heapMem[localMem[2521]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5670;
      end

       5670 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2552]*6 + localMem[2544]] = localMem[2551];
              updateArrayLength(1, localMem[2552], localMem[2544]);
              ip = 5671;
      end

       5671 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2553] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5672;
      end

       5672 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2553]] = localMem[2519];
              ip = 5673;
      end

       5673 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2554] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5674;
      end

       5674 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2554]] = localMem[2519];
              ip = 5675;
      end

       5675 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2555] = localMem[2544] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5676;
      end

       5676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2521]*6 + 0] = localMem[2555];
              updateArrayLength(1, localMem[2521], 0);
              ip = 5677;
      end

       5677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2556] = heapMem[localMem[2521]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5678;
      end

       5678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2556]*6 + localMem[2555]] = localMem[2522];
              updateArrayLength(1, localMem[2556], localMem[2555]);
              ip = 5679;
      end

       5679 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5819;
      end

       5680 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5703;
      end

       5681 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5682;
      end

       5682 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 5683;
      end

       5683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2557] = heapMem[localMem[2521]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5684;
      end

       5684 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2558] = 0; k = arraySizes[localMem[2557]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2557] * NArea + i] == localMem[2514]) localMem[2558] = i + 1;
              end
              ip = 5685;
      end

       5685 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2558] = localMem[2558] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5686;
      end

       5686 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2559] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5687;
      end

       5687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2560] = heapMem[localMem[2559]*6 + localMem[2519]];
              updateArrayLength(2, 0, 0);
              ip = 5688;
      end

       5688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2561] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5689;
      end

       5689 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2562] = heapMem[localMem[2561]*6 + localMem[2519]];
              updateArrayLength(2, 0, 0);
              ip = 5690;
      end

       5690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2563] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5691;
      end

       5691 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2563]] = localMem[2519];
              ip = 5692;
      end

       5692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2564] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5693;
      end

       5693 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2564]] = localMem[2519];
              ip = 5694;
      end

       5694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2565] = heapMem[localMem[2521]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5695;
      end

       5695 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2565] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2558], localMem[2565], arraySizes[localMem[2565]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2558] && i <= arraySizes[localMem[2565]]) begin
                  heapMem[NArea * localMem[2565] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2565] + localMem[2558]] = localMem[2560];                                    // Insert new value
              arraySizes[localMem[2565]] = arraySizes[localMem[2565]] + 1;                              // Increase array size
              ip = 5696;
      end

       5696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2566] = heapMem[localMem[2521]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5697;
      end

       5697 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2566] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2558], localMem[2566], arraySizes[localMem[2566]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2558] && i <= arraySizes[localMem[2566]]) begin
                  heapMem[NArea * localMem[2566] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2566] + localMem[2558]] = localMem[2562];                                    // Insert new value
              arraySizes[localMem[2566]] = arraySizes[localMem[2566]] + 1;                              // Increase array size
              ip = 5698;
      end

       5698 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2567] = heapMem[localMem[2521]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5699;
      end

       5699 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2568] = localMem[2558] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5700;
      end

       5700 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2567] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2568], localMem[2567], arraySizes[localMem[2567]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2568] && i <= arraySizes[localMem[2567]]) begin
                  heapMem[NArea * localMem[2567] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2567] + localMem[2568]] = localMem[2522];                                    // Insert new value
              arraySizes[localMem[2567]] = arraySizes[localMem[2567]] + 1;                              // Increase array size
              ip = 5701;
      end

       5701 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2521]*6 + 0] = heapMem[localMem[2521]*6 + 0] + 1;
              updateArrayLength(1, localMem[2521], 0);
              ip = 5702;
      end

       5702 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5819;
      end

       5703 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5704;
      end

       5704 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5705;
      end

       5705 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2569] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2569] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2569]] = 0;
              ip = 5706;
      end

       5706 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 0] = localMem[2519];
              updateArrayLength(1, localMem[2569], 0);
              ip = 5707;
      end

       5707 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 2] = 0;
              updateArrayLength(1, localMem[2569], 2);
              ip = 5708;
      end

       5708 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2570] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2570] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2570]] = 0;
              ip = 5709;
      end

       5709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 4] = localMem[2570];
              updateArrayLength(1, localMem[2569], 4);
              ip = 5710;
      end

       5710 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2571] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2571] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2571]] = 0;
              ip = 5711;
      end

       5711 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 5] = localMem[2571];
              updateArrayLength(1, localMem[2569], 5);
              ip = 5712;
      end

       5712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 6] = 0;
              updateArrayLength(1, localMem[2569], 6);
              ip = 5713;
      end

       5713 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 3] = localMem[2517];
              updateArrayLength(1, localMem[2569], 3);
              ip = 5714;
      end

       5714 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2517]*6 + 1] = heapMem[localMem[2517]*6 + 1] + 1;
              updateArrayLength(1, localMem[2517], 1);
              ip = 5715;
      end

       5715 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 1] = heapMem[localMem[2517]*6 + 1];
              updateArrayLength(1, localMem[2569], 1);
              ip = 5716;
      end

       5716 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2572] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2572] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2572]] = 0;
              ip = 5717;
      end

       5717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 0] = localMem[2519];
              updateArrayLength(1, localMem[2572], 0);
              ip = 5718;
      end

       5718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 2] = 0;
              updateArrayLength(1, localMem[2572], 2);
              ip = 5719;
      end

       5719 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2573] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2573] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2573]] = 0;
              ip = 5720;
      end

       5720 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 4] = localMem[2573];
              updateArrayLength(1, localMem[2572], 4);
              ip = 5721;
      end

       5721 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2574] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2574] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2574]] = 0;
              ip = 5722;
      end

       5722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 5] = localMem[2574];
              updateArrayLength(1, localMem[2572], 5);
              ip = 5723;
      end

       5723 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 6] = 0;
              updateArrayLength(1, localMem[2572], 6);
              ip = 5724;
      end

       5724 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 3] = localMem[2517];
              updateArrayLength(1, localMem[2572], 3);
              ip = 5725;
      end

       5725 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2517]*6 + 1] = heapMem[localMem[2517]*6 + 1] + 1;
              updateArrayLength(1, localMem[2517], 1);
              ip = 5726;
      end

       5726 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 1] = heapMem[localMem[2517]*6 + 1];
              updateArrayLength(1, localMem[2572], 1);
              ip = 5727;
      end

       5727 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2575] = !heapMem[localMem[2514]*6 + 6];
              ip = 5728;
      end

       5728 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2575] != 0 ? 5780 : 5729;
      end

       5729 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2576] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2576] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2576]] = 0;
              ip = 5730;
      end

       5730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 6] = localMem[2576];
              updateArrayLength(1, localMem[2569], 6);
              ip = 5731;
      end

       5731 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2577] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2577] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2577]] = 0;
              ip = 5732;
      end

       5732 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 6] = localMem[2577];
              updateArrayLength(1, localMem[2572], 6);
              ip = 5733;
      end

       5733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2578] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5734;
      end

       5734 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2579] = heapMem[localMem[2569]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5735;
      end

       5735 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2579] + 0 + i] = heapMem[NArea * localMem[2578] + 0 + i];
                  updateArrayLength(1, localMem[2579], 0 + i);
                end
              end
              ip = 5736;
      end

       5736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2580] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5737;
      end

       5737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2581] = heapMem[localMem[2569]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5738;
      end

       5738 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2581] + 0 + i] = heapMem[NArea * localMem[2580] + 0 + i];
                  updateArrayLength(1, localMem[2581], 0 + i);
                end
              end
              ip = 5739;
      end

       5739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2582] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5740;
      end

       5740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2583] = heapMem[localMem[2569]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5741;
      end

       5741 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2584] = localMem[2519] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5742;
      end

       5742 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2584]) begin
                  heapMem[NArea * localMem[2583] + 0 + i] = heapMem[NArea * localMem[2582] + 0 + i];
                  updateArrayLength(1, localMem[2583], 0 + i);
                end
              end
              ip = 5743;
      end

       5743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2585] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5744;
      end

       5744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2586] = heapMem[localMem[2572]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5745;
      end

       5745 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2586] + 0 + i] = heapMem[NArea * localMem[2585] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2586], 0 + i);
                end
              end
              ip = 5746;
      end

       5746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2587] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5747;
      end

       5747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2588] = heapMem[localMem[2572]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5748;
      end

       5748 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2588] + 0 + i] = heapMem[NArea * localMem[2587] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2588], 0 + i);
                end
              end
              ip = 5749;
      end

       5749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2589] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5750;
      end

       5750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2590] = heapMem[localMem[2572]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5751;
      end

       5751 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2591] = localMem[2519] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5752;
      end

       5752 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2591]) begin
                  heapMem[NArea * localMem[2590] + 0 + i] = heapMem[NArea * localMem[2589] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2590], 0 + i);
                end
              end
              ip = 5753;
      end

       5753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2592] = heapMem[localMem[2569]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5754;
      end

       5754 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2593] = localMem[2592] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5755;
      end

       5755 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2594] = heapMem[localMem[2569]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5756;
      end

       5756 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5757;
      end

       5757 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2595] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5758;
      end

       5758 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5759;
      end

       5759 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2595] >= localMem[2593] ? 5765 : 5760;
      end

       5760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2596] = heapMem[localMem[2594]*6 + localMem[2595]];
              updateArrayLength(2, 0, 0);
              ip = 5761;
      end

       5761 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2596]*6 + 2] = localMem[2569];
              updateArrayLength(1, localMem[2596], 2);
              ip = 5762;
      end

       5762 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5763;
      end

       5763 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2595] = localMem[2595] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5764;
      end

       5764 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5758;
      end

       5765 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5766;
      end

       5766 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2597] = heapMem[localMem[2572]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5767;
      end

       5767 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2598] = localMem[2597] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5768;
      end

       5768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2599] = heapMem[localMem[2572]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5769;
      end

       5769 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5770;
      end

       5770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2600] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5771;
      end

       5771 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5772;
      end

       5772 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2600] >= localMem[2598] ? 5778 : 5773;
      end

       5773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2601] = heapMem[localMem[2599]*6 + localMem[2600]];
              updateArrayLength(2, 0, 0);
              ip = 5774;
      end

       5774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2601]*6 + 2] = localMem[2572];
              updateArrayLength(1, localMem[2601], 2);
              ip = 5775;
      end

       5775 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5776;
      end

       5776 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2600] = localMem[2600] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5777;
      end

       5777 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5771;
      end

       5778 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5779;
      end

       5779 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5795;
      end

       5780 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5781;
      end

       5781 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2602] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2602] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2602]] = 0;
              ip = 5782;
      end

       5782 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2514]*6 + 6] = localMem[2602];
              updateArrayLength(1, localMem[2514], 6);
              ip = 5783;
      end

       5783 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2603] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5784;
      end

       5784 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2604] = heapMem[localMem[2569]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5785;
      end

       5785 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2604] + 0 + i] = heapMem[NArea * localMem[2603] + 0 + i];
                  updateArrayLength(1, localMem[2604], 0 + i);
                end
              end
              ip = 5786;
      end

       5786 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2605] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5787;
      end

       5787 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2606] = heapMem[localMem[2569]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5788;
      end

       5788 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2606] + 0 + i] = heapMem[NArea * localMem[2605] + 0 + i];
                  updateArrayLength(1, localMem[2606], 0 + i);
                end
              end
              ip = 5789;
      end

       5789 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2607] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5790;
      end

       5790 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2608] = heapMem[localMem[2572]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5791;
      end

       5791 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2608] + 0 + i] = heapMem[NArea * localMem[2607] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2608], 0 + i);
                end
              end
              ip = 5792;
      end

       5792 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2609] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5793;
      end

       5793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2610] = heapMem[localMem[2572]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5794;
      end

       5794 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2519]) begin
                  heapMem[NArea * localMem[2610] + 0 + i] = heapMem[NArea * localMem[2609] + localMem[2520] + i];
                  updateArrayLength(1, localMem[2610], 0 + i);
                end
              end
              ip = 5795;
      end

       5795 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5796;
      end

       5796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2569]*6 + 2] = localMem[2514];
              updateArrayLength(1, localMem[2569], 2);
              ip = 5797;
      end

       5797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2572]*6 + 2] = localMem[2514];
              updateArrayLength(1, localMem[2572], 2);
              ip = 5798;
      end

       5798 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2611] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5799;
      end

       5799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2612] = heapMem[localMem[2611]*6 + localMem[2519]];
              updateArrayLength(2, 0, 0);
              ip = 5800;
      end

       5800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2613] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5801;
      end

       5801 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2614] = heapMem[localMem[2613]*6 + localMem[2519]];
              updateArrayLength(2, 0, 0);
              ip = 5802;
      end

       5802 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2615] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5803;
      end

       5803 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2615]*6 + 0] = localMem[2612];
              updateArrayLength(1, localMem[2615], 0);
              ip = 5804;
      end

       5804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2616] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5805;
      end

       5805 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2616]*6 + 0] = localMem[2614];
              updateArrayLength(1, localMem[2616], 0);
              ip = 5806;
      end

       5806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2617] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5807;
      end

       5807 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2617]*6 + 0] = localMem[2569];
              updateArrayLength(1, localMem[2617], 0);
              ip = 5808;
      end

       5808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2618] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5809;
      end

       5809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2618]*6 + 1] = localMem[2572];
              updateArrayLength(1, localMem[2618], 1);
              ip = 5810;
      end

       5810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2514]*6 + 0] = 1;
              updateArrayLength(1, localMem[2514], 0);
              ip = 5811;
      end

       5811 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2619] = heapMem[localMem[2514]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5812;
      end

       5812 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2619]] = 1;
              ip = 5813;
      end

       5813 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2620] = heapMem[localMem[2514]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5814;
      end

       5814 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2620]] = 1;
              ip = 5815;
      end

       5815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2621] = heapMem[localMem[2514]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5816;
      end

       5816 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2621]] = 2;
              ip = 5817;
      end

       5817 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5819;
      end

       5818 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5824;
      end

       5819 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5820;
      end

       5820 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2515] = 1;
              updateArrayLength(2, 0, 0);
              ip = 5821;
      end

       5821 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5824;
      end

       5822 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5823;
      end

       5823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2515] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5824;
      end

       5824 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5825;
      end

       5825 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2515] != 0 ? 5827 : 5826;
      end

       5826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2399] = localMem[2514];
              updateArrayLength(2, 0, 0);
              ip = 5827;
      end

       5827 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5828;
      end

       5828 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6078;
      end

       5829 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5830;
      end

       5830 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2622] = heapMem[localMem[2399]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5831;
      end

       5831 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2623] = 0; k = arraySizes[localMem[2622]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2622] * NArea + i] == 6) localMem[2623] = i + 1;
              end
              ip = 5832;
      end

       5832 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2623] == 0 ? 5837 : 5833;
      end

       5833 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 0] = localMem[2399];
              updateArrayLength(1, localMem[2376], 0);
              ip = 5834;
      end

       5834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 1] = 1;
              updateArrayLength(1, localMem[2376], 1);
              ip = 5835;
      end

       5835 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[2376]*6 + 2] = localMem[2623] - 1;
              updateArrayLength(1, localMem[2376], 2);
              ip = 5836;
      end

       5836 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6085;
      end

       5837 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5838;
      end

       5838 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
              j = 0; k = arraySizes[localMem[2622]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2622] * NArea + i] < 6) j = j + 1;
              end
              localMem[2624] = j;
              ip = 5839;
      end

       5839 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2625] = !heapMem[localMem[2399]*6 + 6];
              ip = 5840;
      end

       5840 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2625] == 0 ? 5845 : 5841;
      end

       5841 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 0] = localMem[2399];
              updateArrayLength(1, localMem[2376], 0);
              ip = 5842;
      end

       5842 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 1] = 0;
              updateArrayLength(1, localMem[2376], 1);
              ip = 5843;
      end

       5843 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*6 + 2] = localMem[2624];
              updateArrayLength(1, localMem[2376], 2);
              ip = 5844;
      end

       5844 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6085;
      end

       5845 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5846;
      end

       5846 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2626] = heapMem[localMem[2399]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5847;
      end

       5847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2627] = heapMem[localMem[2626]*6 + localMem[2624]];
              updateArrayLength(2, 0, 0);
              ip = 5848;
      end

       5848 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5849;
      end

       5849 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2629] = heapMem[localMem[2627]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5850;
      end

       5850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2630] = heapMem[localMem[2627]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5851;
      end

       5851 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2631] = heapMem[localMem[2630]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5852;
      end

       5852 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2629] <  localMem[2631] ? 6072 : 5853;
      end

       5853 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2632] = localMem[2631];
              updateArrayLength(2, 0, 0);
              ip = 5854;
      end

       5854 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2632] = localMem[2632] >> 1;
              ip = 5855;
      end

       5855 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2633] = localMem[2632] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5856;
      end

       5856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2634] = heapMem[localMem[2627]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5857;
      end

       5857 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2634] == 0 ? 5954 : 5858;
      end

       5858 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2635] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2635] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2635]] = 0;
              ip = 5859;
      end

       5859 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 0] = localMem[2632];
              updateArrayLength(1, localMem[2635], 0);
              ip = 5860;
      end

       5860 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 2] = 0;
              updateArrayLength(1, localMem[2635], 2);
              ip = 5861;
      end

       5861 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2636] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2636] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2636]] = 0;
              ip = 5862;
      end

       5862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 4] = localMem[2636];
              updateArrayLength(1, localMem[2635], 4);
              ip = 5863;
      end

       5863 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2637] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2637] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2637]] = 0;
              ip = 5864;
      end

       5864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 5] = localMem[2637];
              updateArrayLength(1, localMem[2635], 5);
              ip = 5865;
      end

       5865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 6] = 0;
              updateArrayLength(1, localMem[2635], 6);
              ip = 5866;
      end

       5866 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 3] = localMem[2630];
              updateArrayLength(1, localMem[2635], 3);
              ip = 5867;
      end

       5867 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2630]*6 + 1] = heapMem[localMem[2630]*6 + 1] + 1;
              updateArrayLength(1, localMem[2630], 1);
              ip = 5868;
      end

       5868 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 1] = heapMem[localMem[2630]*6 + 1];
              updateArrayLength(1, localMem[2635], 1);
              ip = 5869;
      end

       5869 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2638] = !heapMem[localMem[2627]*6 + 6];
              ip = 5870;
      end

       5870 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2638] != 0 ? 5899 : 5871;
      end

       5871 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2639] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2639] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2639]] = 0;
              ip = 5872;
      end

       5872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 6] = localMem[2639];
              updateArrayLength(1, localMem[2635], 6);
              ip = 5873;
      end

       5873 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2640] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5874;
      end

       5874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2641] = heapMem[localMem[2635]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5875;
      end

       5875 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2641] + 0 + i] = heapMem[NArea * localMem[2640] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2641], 0 + i);
                end
              end
              ip = 5876;
      end

       5876 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2642] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5877;
      end

       5877 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2643] = heapMem[localMem[2635]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5878;
      end

       5878 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2643] + 0 + i] = heapMem[NArea * localMem[2642] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2643], 0 + i);
                end
              end
              ip = 5879;
      end

       5879 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2644] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5880;
      end

       5880 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2645] = heapMem[localMem[2635]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5881;
      end

       5881 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2646] = localMem[2632] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5882;
      end

       5882 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2646]) begin
                  heapMem[NArea * localMem[2645] + 0 + i] = heapMem[NArea * localMem[2644] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2645], 0 + i);
                end
              end
              ip = 5883;
      end

       5883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2647] = heapMem[localMem[2635]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5884;
      end

       5884 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2648] = localMem[2647] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5885;
      end

       5885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2649] = heapMem[localMem[2635]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5886;
      end

       5886 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5887;
      end

       5887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2650] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5888;
      end

       5888 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5889;
      end

       5889 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2650] >= localMem[2648] ? 5895 : 5890;
      end

       5890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2651] = heapMem[localMem[2649]*6 + localMem[2650]];
              updateArrayLength(2, 0, 0);
              ip = 5891;
      end

       5891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2651]*6 + 2] = localMem[2635];
              updateArrayLength(1, localMem[2651], 2);
              ip = 5892;
      end

       5892 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5893;
      end

       5893 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2650] = localMem[2650] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5894;
      end

       5894 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5888;
      end

       5895 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5896;
      end

       5896 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2652] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5897;
      end

       5897 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2652]] = localMem[2633];
              ip = 5898;
      end

       5898 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5906;
      end

       5899 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5900;
      end

       5900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2653] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5901;
      end

       5901 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2654] = heapMem[localMem[2635]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5902;
      end

       5902 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2654] + 0 + i] = heapMem[NArea * localMem[2653] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2654], 0 + i);
                end
              end
              ip = 5903;
      end

       5903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2655] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5904;
      end

       5904 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2656] = heapMem[localMem[2635]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5905;
      end

       5905 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2656] + 0 + i] = heapMem[NArea * localMem[2655] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2656], 0 + i);
                end
              end
              ip = 5906;
      end

       5906 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5907;
      end

       5907 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2627]*6 + 0] = localMem[2632];
              updateArrayLength(1, localMem[2627], 0);
              ip = 5908;
      end

       5908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2635]*6 + 2] = localMem[2634];
              updateArrayLength(1, localMem[2635], 2);
              ip = 5909;
      end

       5909 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2657] = heapMem[localMem[2634]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5910;
      end

       5910 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2658] = heapMem[localMem[2634]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5911;
      end

       5911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2659] = heapMem[localMem[2658]*6 + localMem[2657]];
              updateArrayLength(2, 0, 0);
              ip = 5912;
      end

       5912 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2659] != localMem[2627] ? 5931 : 5913;
      end

       5913 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2660] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5914;
      end

       5914 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2661] = heapMem[localMem[2660]*6 + localMem[2632]];
              updateArrayLength(2, 0, 0);
              ip = 5915;
      end

       5915 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2662] = heapMem[localMem[2634]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5916;
      end

       5916 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2662]*6 + localMem[2657]] = localMem[2661];
              updateArrayLength(1, localMem[2662], localMem[2657]);
              ip = 5917;
      end

       5917 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2663] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5918;
      end

       5918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2664] = heapMem[localMem[2663]*6 + localMem[2632]];
              updateArrayLength(2, 0, 0);
              ip = 5919;
      end

       5919 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2665] = heapMem[localMem[2634]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5920;
      end

       5920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2665]*6 + localMem[2657]] = localMem[2664];
              updateArrayLength(1, localMem[2665], localMem[2657]);
              ip = 5921;
      end

       5921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2666] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5922;
      end

       5922 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2666]] = localMem[2632];
              ip = 5923;
      end

       5923 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2667] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5924;
      end

       5924 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2667]] = localMem[2632];
              ip = 5925;
      end

       5925 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2668] = localMem[2657] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5926;
      end

       5926 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2634]*6 + 0] = localMem[2668];
              updateArrayLength(1, localMem[2634], 0);
              ip = 5927;
      end

       5927 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2669] = heapMem[localMem[2634]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5928;
      end

       5928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2669]*6 + localMem[2668]] = localMem[2635];
              updateArrayLength(1, localMem[2669], localMem[2668]);
              ip = 5929;
      end

       5929 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6069;
      end

       5930 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5953;
      end

       5931 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5932;
      end

       5932 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 5933;
      end

       5933 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2670] = heapMem[localMem[2634]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5934;
      end

       5934 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2671] = 0; k = arraySizes[localMem[2670]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2670] * NArea + i] == localMem[2627]) localMem[2671] = i + 1;
              end
              ip = 5935;
      end

       5935 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2671] = localMem[2671] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5936;
      end

       5936 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2672] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5937;
      end

       5937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2673] = heapMem[localMem[2672]*6 + localMem[2632]];
              updateArrayLength(2, 0, 0);
              ip = 5938;
      end

       5938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2674] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5939;
      end

       5939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2675] = heapMem[localMem[2674]*6 + localMem[2632]];
              updateArrayLength(2, 0, 0);
              ip = 5940;
      end

       5940 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2676] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5941;
      end

       5941 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2676]] = localMem[2632];
              ip = 5942;
      end

       5942 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2677] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5943;
      end

       5943 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2677]] = localMem[2632];
              ip = 5944;
      end

       5944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2678] = heapMem[localMem[2634]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5945;
      end

       5945 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2678] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2671], localMem[2678], arraySizes[localMem[2678]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2671] && i <= arraySizes[localMem[2678]]) begin
                  heapMem[NArea * localMem[2678] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2678] + localMem[2671]] = localMem[2673];                                    // Insert new value
              arraySizes[localMem[2678]] = arraySizes[localMem[2678]] + 1;                              // Increase array size
              ip = 5946;
      end

       5946 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2679] = heapMem[localMem[2634]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5947;
      end

       5947 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2679] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2671], localMem[2679], arraySizes[localMem[2679]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2671] && i <= arraySizes[localMem[2679]]) begin
                  heapMem[NArea * localMem[2679] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2679] + localMem[2671]] = localMem[2675];                                    // Insert new value
              arraySizes[localMem[2679]] = arraySizes[localMem[2679]] + 1;                              // Increase array size
              ip = 5948;
      end

       5948 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2680] = heapMem[localMem[2634]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5949;
      end

       5949 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2681] = localMem[2671] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5950;
      end

       5950 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2680] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2681], localMem[2680], arraySizes[localMem[2680]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2681] && i <= arraySizes[localMem[2680]]) begin
                  heapMem[NArea * localMem[2680] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2680] + localMem[2681]] = localMem[2635];                                    // Insert new value
              arraySizes[localMem[2680]] = arraySizes[localMem[2680]] + 1;                              // Increase array size
              ip = 5951;
      end

       5951 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2634]*6 + 0] = heapMem[localMem[2634]*6 + 0] + 1;
              updateArrayLength(1, localMem[2634], 0);
              ip = 5952;
      end

       5952 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6069;
      end

       5953 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5954;
      end

       5954 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5955;
      end

       5955 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2682] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2682] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2682]] = 0;
              ip = 5956;
      end

       5956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 0] = localMem[2632];
              updateArrayLength(1, localMem[2682], 0);
              ip = 5957;
      end

       5957 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 2] = 0;
              updateArrayLength(1, localMem[2682], 2);
              ip = 5958;
      end

       5958 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2683] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2683] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2683]] = 0;
              ip = 5959;
      end

       5959 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 4] = localMem[2683];
              updateArrayLength(1, localMem[2682], 4);
              ip = 5960;
      end

       5960 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2684] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2684] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2684]] = 0;
              ip = 5961;
      end

       5961 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 5] = localMem[2684];
              updateArrayLength(1, localMem[2682], 5);
              ip = 5962;
      end

       5962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 6] = 0;
              updateArrayLength(1, localMem[2682], 6);
              ip = 5963;
      end

       5963 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 3] = localMem[2630];
              updateArrayLength(1, localMem[2682], 3);
              ip = 5964;
      end

       5964 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2630]*6 + 1] = heapMem[localMem[2630]*6 + 1] + 1;
              updateArrayLength(1, localMem[2630], 1);
              ip = 5965;
      end

       5965 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 1] = heapMem[localMem[2630]*6 + 1];
              updateArrayLength(1, localMem[2682], 1);
              ip = 5966;
      end

       5966 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2685] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2685] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2685]] = 0;
              ip = 5967;
      end

       5967 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 0] = localMem[2632];
              updateArrayLength(1, localMem[2685], 0);
              ip = 5968;
      end

       5968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 2] = 0;
              updateArrayLength(1, localMem[2685], 2);
              ip = 5969;
      end

       5969 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2686] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2686] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2686]] = 0;
              ip = 5970;
      end

       5970 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 4] = localMem[2686];
              updateArrayLength(1, localMem[2685], 4);
              ip = 5971;
      end

       5971 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2687] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2687] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2687]] = 0;
              ip = 5972;
      end

       5972 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 5] = localMem[2687];
              updateArrayLength(1, localMem[2685], 5);
              ip = 5973;
      end

       5973 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 6] = 0;
              updateArrayLength(1, localMem[2685], 6);
              ip = 5974;
      end

       5974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 3] = localMem[2630];
              updateArrayLength(1, localMem[2685], 3);
              ip = 5975;
      end

       5975 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2630]*6 + 1] = heapMem[localMem[2630]*6 + 1] + 1;
              updateArrayLength(1, localMem[2630], 1);
              ip = 5976;
      end

       5976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 1] = heapMem[localMem[2630]*6 + 1];
              updateArrayLength(1, localMem[2685], 1);
              ip = 5977;
      end

       5977 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2688] = !heapMem[localMem[2627]*6 + 6];
              ip = 5978;
      end

       5978 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2688] != 0 ? 6030 : 5979;
      end

       5979 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2689] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2689] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2689]] = 0;
              ip = 5980;
      end

       5980 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 6] = localMem[2689];
              updateArrayLength(1, localMem[2682], 6);
              ip = 5981;
      end

       5981 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2690] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2690] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2690]] = 0;
              ip = 5982;
      end

       5982 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 6] = localMem[2690];
              updateArrayLength(1, localMem[2685], 6);
              ip = 5983;
      end

       5983 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2691] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5984;
      end

       5984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2692] = heapMem[localMem[2682]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5985;
      end

       5985 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2692] + 0 + i] = heapMem[NArea * localMem[2691] + 0 + i];
                  updateArrayLength(1, localMem[2692], 0 + i);
                end
              end
              ip = 5986;
      end

       5986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2693] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5987;
      end

       5987 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2694] = heapMem[localMem[2682]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5988;
      end

       5988 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2694] + 0 + i] = heapMem[NArea * localMem[2693] + 0 + i];
                  updateArrayLength(1, localMem[2694], 0 + i);
                end
              end
              ip = 5989;
      end

       5989 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2695] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5990;
      end

       5990 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2696] = heapMem[localMem[2682]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5991;
      end

       5991 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2697] = localMem[2632] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5992;
      end

       5992 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2697]) begin
                  heapMem[NArea * localMem[2696] + 0 + i] = heapMem[NArea * localMem[2695] + 0 + i];
                  updateArrayLength(1, localMem[2696], 0 + i);
                end
              end
              ip = 5993;
      end

       5993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2698] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5994;
      end

       5994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2699] = heapMem[localMem[2685]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5995;
      end

       5995 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2699] + 0 + i] = heapMem[NArea * localMem[2698] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2699], 0 + i);
                end
              end
              ip = 5996;
      end

       5996 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2700] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5997;
      end

       5997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2701] = heapMem[localMem[2685]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5998;
      end

       5998 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2701] + 0 + i] = heapMem[NArea * localMem[2700] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2701], 0 + i);
                end
              end
              ip = 5999;
      end

       5999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2702] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6000;
      end

       6000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2703] = heapMem[localMem[2685]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6001;
      end

       6001 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2704] = localMem[2632] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6002;
      end

       6002 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2704]) begin
                  heapMem[NArea * localMem[2703] + 0 + i] = heapMem[NArea * localMem[2702] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2703], 0 + i);
                end
              end
              ip = 6003;
      end

       6003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2705] = heapMem[localMem[2682]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6004;
      end

       6004 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2706] = localMem[2705] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6005;
      end

       6005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2707] = heapMem[localMem[2682]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6006;
      end

       6006 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6007;
      end

       6007 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2708] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6008;
      end

       6008 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6009;
      end

       6009 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2708] >= localMem[2706] ? 6015 : 6010;
      end

       6010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2709] = heapMem[localMem[2707]*6 + localMem[2708]];
              updateArrayLength(2, 0, 0);
              ip = 6011;
      end

       6011 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2709]*6 + 2] = localMem[2682];
              updateArrayLength(1, localMem[2709], 2);
              ip = 6012;
      end

       6012 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6013;
      end

       6013 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2708] = localMem[2708] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6014;
      end

       6014 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6008;
      end

       6015 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6016;
      end

       6016 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2710] = heapMem[localMem[2685]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6017;
      end

       6017 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2711] = localMem[2710] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6018;
      end

       6018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2712] = heapMem[localMem[2685]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6019;
      end

       6019 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6020;
      end

       6020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2713] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6021;
      end

       6021 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6022;
      end

       6022 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2713] >= localMem[2711] ? 6028 : 6023;
      end

       6023 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2714] = heapMem[localMem[2712]*6 + localMem[2713]];
              updateArrayLength(2, 0, 0);
              ip = 6024;
      end

       6024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2714]*6 + 2] = localMem[2685];
              updateArrayLength(1, localMem[2714], 2);
              ip = 6025;
      end

       6025 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6026;
      end

       6026 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2713] = localMem[2713] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6027;
      end

       6027 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6021;
      end

       6028 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6029;
      end

       6029 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6045;
      end

       6030 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6031;
      end

       6031 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2715] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2715] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2715]] = 0;
              ip = 6032;
      end

       6032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2627]*6 + 6] = localMem[2715];
              updateArrayLength(1, localMem[2627], 6);
              ip = 6033;
      end

       6033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2716] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6034;
      end

       6034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2717] = heapMem[localMem[2682]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6035;
      end

       6035 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2717] + 0 + i] = heapMem[NArea * localMem[2716] + 0 + i];
                  updateArrayLength(1, localMem[2717], 0 + i);
                end
              end
              ip = 6036;
      end

       6036 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2718] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6037;
      end

       6037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2719] = heapMem[localMem[2682]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6038;
      end

       6038 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2719] + 0 + i] = heapMem[NArea * localMem[2718] + 0 + i];
                  updateArrayLength(1, localMem[2719], 0 + i);
                end
              end
              ip = 6039;
      end

       6039 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2720] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6040;
      end

       6040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2721] = heapMem[localMem[2685]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6041;
      end

       6041 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2721] + 0 + i] = heapMem[NArea * localMem[2720] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2721], 0 + i);
                end
              end
              ip = 6042;
      end

       6042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2722] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6043;
      end

       6043 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2723] = heapMem[localMem[2685]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6044;
      end

       6044 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2632]) begin
                  heapMem[NArea * localMem[2723] + 0 + i] = heapMem[NArea * localMem[2722] + localMem[2633] + i];
                  updateArrayLength(1, localMem[2723], 0 + i);
                end
              end
              ip = 6045;
      end

       6045 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6046;
      end

       6046 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2682]*6 + 2] = localMem[2627];
              updateArrayLength(1, localMem[2682], 2);
              ip = 6047;
      end

       6047 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2685]*6 + 2] = localMem[2627];
              updateArrayLength(1, localMem[2685], 2);
              ip = 6048;
      end

       6048 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2724] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6049;
      end

       6049 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2725] = heapMem[localMem[2724]*6 + localMem[2632]];
              updateArrayLength(2, 0, 0);
              ip = 6050;
      end

       6050 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2726] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6051;
      end

       6051 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2727] = heapMem[localMem[2726]*6 + localMem[2632]];
              updateArrayLength(2, 0, 0);
              ip = 6052;
      end

       6052 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2728] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6053;
      end

       6053 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2728]*6 + 0] = localMem[2725];
              updateArrayLength(1, localMem[2728], 0);
              ip = 6054;
      end

       6054 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2729] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6055;
      end

       6055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2729]*6 + 0] = localMem[2727];
              updateArrayLength(1, localMem[2729], 0);
              ip = 6056;
      end

       6056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2730] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6057;
      end

       6057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2730]*6 + 0] = localMem[2682];
              updateArrayLength(1, localMem[2730], 0);
              ip = 6058;
      end

       6058 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2731] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6059;
      end

       6059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2731]*6 + 1] = localMem[2685];
              updateArrayLength(1, localMem[2731], 1);
              ip = 6060;
      end

       6060 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2627]*6 + 0] = 1;
              updateArrayLength(1, localMem[2627], 0);
              ip = 6061;
      end

       6061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2732] = heapMem[localMem[2627]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6062;
      end

       6062 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2732]] = 1;
              ip = 6063;
      end

       6063 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2733] = heapMem[localMem[2627]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6064;
      end

       6064 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2733]] = 1;
              ip = 6065;
      end

       6065 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2734] = heapMem[localMem[2627]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6066;
      end

       6066 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2734]] = 2;
              ip = 6067;
      end

       6067 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6069;
      end

       6068 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6074;
      end

       6069 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6070;
      end

       6070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2628] = 1;
              updateArrayLength(2, 0, 0);
              ip = 6071;
      end

       6071 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6074;
      end

       6072 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6073;
      end

       6073 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2628] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6074;
      end

       6074 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6075;
      end

       6075 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2628] != 0 ? 6077 : 6076;
      end

       6076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2399] = localMem[2627];
              updateArrayLength(2, 0, 0);
              ip = 6077;
      end

       6077 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6078;
      end

       6078 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6079;
      end

       6079 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2507] = localMem[2507] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6080;
      end

       6080 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5582;
      end

       6081 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6082;
      end

       6082 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
            ip = 6083;
      end

       6083 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6084;
      end

       6084 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6085;
      end

       6085 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6086;
      end

       6086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2735] = heapMem[localMem[2376]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6087;
      end

       6087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2736] = heapMem[localMem[2376]*6 + 1];
              updateArrayLength(2, 0, 0);
              ip = 6088;
      end

       6088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2737] = heapMem[localMem[2376]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 6089;
      end

       6089 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2736] != 1 ? 6093 : 6090;
      end

       6090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2738] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6091;
      end

       6091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2738]*6 + localMem[2737]] = 66;
              updateArrayLength(1, localMem[2738], localMem[2737]);
              ip = 6092;
      end

       6092 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6339;
      end

       6093 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6094;
      end

       6094 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2736] != 2 ? 6102 : 6095;
      end

       6095 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2739] = localMem[2737] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6096;
      end

       6096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2740] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6097;
      end

       6097 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2740] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2739], localMem[2740], arraySizes[localMem[2740]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2739] && i <= arraySizes[localMem[2740]]) begin
                  heapMem[NArea * localMem[2740] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2740] + localMem[2739]] = 6;                                    // Insert new value
              arraySizes[localMem[2740]] = arraySizes[localMem[2740]] + 1;                              // Increase array size
              ip = 6098;
      end

       6098 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2741] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6099;
      end

       6099 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2741] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2739], localMem[2741], arraySizes[localMem[2741]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2739] && i <= arraySizes[localMem[2741]]) begin
                  heapMem[NArea * localMem[2741] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2741] + localMem[2739]] = 66;                                    // Insert new value
              arraySizes[localMem[2741]] = arraySizes[localMem[2741]] + 1;                              // Increase array size
              ip = 6100;
      end

       6100 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2735]*6 + 0] = heapMem[localMem[2735]*6 + 0] + 1;
              updateArrayLength(1, localMem[2735], 0);
              ip = 6101;
      end

       6101 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6108;
      end

       6102 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6103;
      end

       6103 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2742] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6104;
      end

       6104 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2742] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2737], localMem[2742], arraySizes[localMem[2742]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2737] && i <= arraySizes[localMem[2742]]) begin
                  heapMem[NArea * localMem[2742] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2742] + localMem[2737]] = 6;                                    // Insert new value
              arraySizes[localMem[2742]] = arraySizes[localMem[2742]] + 1;                              // Increase array size
              ip = 6105;
      end

       6105 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2743] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6106;
      end

       6106 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2743] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2737], localMem[2743], arraySizes[localMem[2743]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2737] && i <= arraySizes[localMem[2743]]) begin
                  heapMem[NArea * localMem[2743] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2743] + localMem[2737]] = 66;                                    // Insert new value
              arraySizes[localMem[2743]] = arraySizes[localMem[2743]] + 1;                              // Increase array size
              ip = 6107;
      end

       6107 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2735]*6 + 0] = heapMem[localMem[2735]*6 + 0] + 1;
              updateArrayLength(1, localMem[2735], 0);
              ip = 6108;
      end

       6108 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6109;
      end

       6109 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*6 + 0] = heapMem[localMem[0]*6 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 6110;
      end

       6110 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6111;
      end

       6111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2745] = heapMem[localMem[2735]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6112;
      end

       6112 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2746] = heapMem[localMem[2735]*6 + 3];
              updateArrayLength(2, 0, 0);
              ip = 6113;
      end

       6113 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2747] = heapMem[localMem[2746]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 6114;
      end

       6114 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2745] <  localMem[2747] ? 6334 : 6115;
      end

       6115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2748] = localMem[2747];
              updateArrayLength(2, 0, 0);
              ip = 6116;
      end

       6116 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2748] = localMem[2748] >> 1;
              ip = 6117;
      end

       6117 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2749] = localMem[2748] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6118;
      end

       6118 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2750] = heapMem[localMem[2735]*6 + 2];
              updateArrayLength(2, 0, 0);
              ip = 6119;
      end

       6119 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2750] == 0 ? 6216 : 6120;
      end

       6120 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2751] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2751] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2751]] = 0;
              ip = 6121;
      end

       6121 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 0] = localMem[2748];
              updateArrayLength(1, localMem[2751], 0);
              ip = 6122;
      end

       6122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 2] = 0;
              updateArrayLength(1, localMem[2751], 2);
              ip = 6123;
      end

       6123 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2752] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2752] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2752]] = 0;
              ip = 6124;
      end

       6124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 4] = localMem[2752];
              updateArrayLength(1, localMem[2751], 4);
              ip = 6125;
      end

       6125 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2753] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2753] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2753]] = 0;
              ip = 6126;
      end

       6126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 5] = localMem[2753];
              updateArrayLength(1, localMem[2751], 5);
              ip = 6127;
      end

       6127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 6] = 0;
              updateArrayLength(1, localMem[2751], 6);
              ip = 6128;
      end

       6128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 3] = localMem[2746];
              updateArrayLength(1, localMem[2751], 3);
              ip = 6129;
      end

       6129 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2746]*6 + 1] = heapMem[localMem[2746]*6 + 1] + 1;
              updateArrayLength(1, localMem[2746], 1);
              ip = 6130;
      end

       6130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 1] = heapMem[localMem[2746]*6 + 1];
              updateArrayLength(1, localMem[2751], 1);
              ip = 6131;
      end

       6131 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2754] = !heapMem[localMem[2735]*6 + 6];
              ip = 6132;
      end

       6132 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2754] != 0 ? 6161 : 6133;
      end

       6133 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2755] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2755] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2755]] = 0;
              ip = 6134;
      end

       6134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 6] = localMem[2755];
              updateArrayLength(1, localMem[2751], 6);
              ip = 6135;
      end

       6135 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2756] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6136;
      end

       6136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2757] = heapMem[localMem[2751]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6137;
      end

       6137 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2757] + 0 + i] = heapMem[NArea * localMem[2756] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2757], 0 + i);
                end
              end
              ip = 6138;
      end

       6138 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2758] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6139;
      end

       6139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2759] = heapMem[localMem[2751]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6140;
      end

       6140 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2759] + 0 + i] = heapMem[NArea * localMem[2758] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2759], 0 + i);
                end
              end
              ip = 6141;
      end

       6141 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2760] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6142;
      end

       6142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2761] = heapMem[localMem[2751]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6143;
      end

       6143 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2762] = localMem[2748] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6144;
      end

       6144 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2762]) begin
                  heapMem[NArea * localMem[2761] + 0 + i] = heapMem[NArea * localMem[2760] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2761], 0 + i);
                end
              end
              ip = 6145;
      end

       6145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2763] = heapMem[localMem[2751]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6146;
      end

       6146 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2764] = localMem[2763] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6147;
      end

       6147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2765] = heapMem[localMem[2751]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6148;
      end

       6148 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6149;
      end

       6149 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2766] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6150;
      end

       6150 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6151;
      end

       6151 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2766] >= localMem[2764] ? 6157 : 6152;
      end

       6152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2767] = heapMem[localMem[2765]*6 + localMem[2766]];
              updateArrayLength(2, 0, 0);
              ip = 6153;
      end

       6153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2767]*6 + 2] = localMem[2751];
              updateArrayLength(1, localMem[2767], 2);
              ip = 6154;
      end

       6154 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6155;
      end

       6155 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2766] = localMem[2766] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6156;
      end

       6156 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6150;
      end

       6157 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6158;
      end

       6158 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2768] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6159;
      end

       6159 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2768]] = localMem[2749];
              ip = 6160;
      end

       6160 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6168;
      end

       6161 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6162;
      end

       6162 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2769] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6163;
      end

       6163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2770] = heapMem[localMem[2751]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6164;
      end

       6164 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2770] + 0 + i] = heapMem[NArea * localMem[2769] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2770], 0 + i);
                end
              end
              ip = 6165;
      end

       6165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2771] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6166;
      end

       6166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2772] = heapMem[localMem[2751]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6167;
      end

       6167 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2772] + 0 + i] = heapMem[NArea * localMem[2771] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2772], 0 + i);
                end
              end
              ip = 6168;
      end

       6168 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6169;
      end

       6169 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2735]*6 + 0] = localMem[2748];
              updateArrayLength(1, localMem[2735], 0);
              ip = 6170;
      end

       6170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2751]*6 + 2] = localMem[2750];
              updateArrayLength(1, localMem[2751], 2);
              ip = 6171;
      end

       6171 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2773] = heapMem[localMem[2750]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6172;
      end

       6172 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2774] = heapMem[localMem[2750]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6173;
      end

       6173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2775] = heapMem[localMem[2774]*6 + localMem[2773]];
              updateArrayLength(2, 0, 0);
              ip = 6174;
      end

       6174 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2775] != localMem[2735] ? 6193 : 6175;
      end

       6175 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2776] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6176;
      end

       6176 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2777] = heapMem[localMem[2776]*6 + localMem[2748]];
              updateArrayLength(2, 0, 0);
              ip = 6177;
      end

       6177 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2778] = heapMem[localMem[2750]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6178;
      end

       6178 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2778]*6 + localMem[2773]] = localMem[2777];
              updateArrayLength(1, localMem[2778], localMem[2773]);
              ip = 6179;
      end

       6179 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2779] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6180;
      end

       6180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2780] = heapMem[localMem[2779]*6 + localMem[2748]];
              updateArrayLength(2, 0, 0);
              ip = 6181;
      end

       6181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2781] = heapMem[localMem[2750]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6182;
      end

       6182 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2781]*6 + localMem[2773]] = localMem[2780];
              updateArrayLength(1, localMem[2781], localMem[2773]);
              ip = 6183;
      end

       6183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2782] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6184;
      end

       6184 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2782]] = localMem[2748];
              ip = 6185;
      end

       6185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2783] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6186;
      end

       6186 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2783]] = localMem[2748];
              ip = 6187;
      end

       6187 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2784] = localMem[2773] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6188;
      end

       6188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2750]*6 + 0] = localMem[2784];
              updateArrayLength(1, localMem[2750], 0);
              ip = 6189;
      end

       6189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2785] = heapMem[localMem[2750]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6190;
      end

       6190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2785]*6 + localMem[2784]] = localMem[2751];
              updateArrayLength(1, localMem[2785], localMem[2784]);
              ip = 6191;
      end

       6191 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6331;
      end

       6192 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6215;
      end

       6193 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6194;
      end

       6194 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
            ip = 6195;
      end

       6195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2786] = heapMem[localMem[2750]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6196;
      end

       6196 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[2787] = 0; k = arraySizes[localMem[2786]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[2786] * NArea + i] == localMem[2735]) localMem[2787] = i + 1;
              end
              ip = 6197;
      end

       6197 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2787] = localMem[2787] - 1;
              updateArrayLength(2, 0, 0);
              ip = 6198;
      end

       6198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2788] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6199;
      end

       6199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2789] = heapMem[localMem[2788]*6 + localMem[2748]];
              updateArrayLength(2, 0, 0);
              ip = 6200;
      end

       6200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2790] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6201;
      end

       6201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2791] = heapMem[localMem[2790]*6 + localMem[2748]];
              updateArrayLength(2, 0, 0);
              ip = 6202;
      end

       6202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2792] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6203;
      end

       6203 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2792]] = localMem[2748];
              ip = 6204;
      end

       6204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2793] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6205;
      end

       6205 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2793]] = localMem[2748];
              ip = 6206;
      end

       6206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2794] = heapMem[localMem[2750]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6207;
      end

       6207 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2794] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2787], localMem[2794], arraySizes[localMem[2794]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2787] && i <= arraySizes[localMem[2794]]) begin
                  heapMem[NArea * localMem[2794] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2794] + localMem[2787]] = localMem[2789];                                    // Insert new value
              arraySizes[localMem[2794]] = arraySizes[localMem[2794]] + 1;                              // Increase array size
              ip = 6208;
      end

       6208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2795] = heapMem[localMem[2750]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6209;
      end

       6209 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2795] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2787], localMem[2795], arraySizes[localMem[2795]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2787] && i <= arraySizes[localMem[2795]]) begin
                  heapMem[NArea * localMem[2795] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2795] + localMem[2787]] = localMem[2791];                                    // Insert new value
              arraySizes[localMem[2795]] = arraySizes[localMem[2795]] + 1;                              // Increase array size
              ip = 6210;
      end

       6210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2796] = heapMem[localMem[2750]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6211;
      end

       6211 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2797] = localMem[2787] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6212;
      end

       6212 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2796] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2797], localMem[2796], arraySizes[localMem[2796]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2797] && i <= arraySizes[localMem[2796]]) begin
                  heapMem[NArea * localMem[2796] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2796] + localMem[2797]] = localMem[2751];                                    // Insert new value
              arraySizes[localMem[2796]] = arraySizes[localMem[2796]] + 1;                              // Increase array size
              ip = 6213;
      end

       6213 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2750]*6 + 0] = heapMem[localMem[2750]*6 + 0] + 1;
              updateArrayLength(1, localMem[2750], 0);
              ip = 6214;
      end

       6214 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6331;
      end

       6215 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6216;
      end

       6216 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6217;
      end

       6217 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2798] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2798] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2798]] = 0;
              ip = 6218;
      end

       6218 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 0] = localMem[2748];
              updateArrayLength(1, localMem[2798], 0);
              ip = 6219;
      end

       6219 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 2] = 0;
              updateArrayLength(1, localMem[2798], 2);
              ip = 6220;
      end

       6220 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2799] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2799] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2799]] = 0;
              ip = 6221;
      end

       6221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 4] = localMem[2799];
              updateArrayLength(1, localMem[2798], 4);
              ip = 6222;
      end

       6222 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2800] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2800] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2800]] = 0;
              ip = 6223;
      end

       6223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 5] = localMem[2800];
              updateArrayLength(1, localMem[2798], 5);
              ip = 6224;
      end

       6224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 6] = 0;
              updateArrayLength(1, localMem[2798], 6);
              ip = 6225;
      end

       6225 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 3] = localMem[2746];
              updateArrayLength(1, localMem[2798], 3);
              ip = 6226;
      end

       6226 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2746]*6 + 1] = heapMem[localMem[2746]*6 + 1] + 1;
              updateArrayLength(1, localMem[2746], 1);
              ip = 6227;
      end

       6227 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 1] = heapMem[localMem[2746]*6 + 1];
              updateArrayLength(1, localMem[2798], 1);
              ip = 6228;
      end

       6228 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2801] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2801] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2801]] = 0;
              ip = 6229;
      end

       6229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 0] = localMem[2748];
              updateArrayLength(1, localMem[2801], 0);
              ip = 6230;
      end

       6230 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 2] = 0;
              updateArrayLength(1, localMem[2801], 2);
              ip = 6231;
      end

       6231 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2802] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2802] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2802]] = 0;
              ip = 6232;
      end

       6232 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 4] = localMem[2802];
              updateArrayLength(1, localMem[2801], 4);
              ip = 6233;
      end

       6233 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2803] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2803] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2803]] = 0;
              ip = 6234;
      end

       6234 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 5] = localMem[2803];
              updateArrayLength(1, localMem[2801], 5);
              ip = 6235;
      end

       6235 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 6] = 0;
              updateArrayLength(1, localMem[2801], 6);
              ip = 6236;
      end

       6236 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 3] = localMem[2746];
              updateArrayLength(1, localMem[2801], 3);
              ip = 6237;
      end

       6237 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2746]*6 + 1] = heapMem[localMem[2746]*6 + 1] + 1;
              updateArrayLength(1, localMem[2746], 1);
              ip = 6238;
      end

       6238 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 1] = heapMem[localMem[2746]*6 + 1];
              updateArrayLength(1, localMem[2801], 1);
              ip = 6239;
      end

       6239 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2804] = !heapMem[localMem[2735]*6 + 6];
              ip = 6240;
      end

       6240 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2804] != 0 ? 6292 : 6241;
      end

       6241 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2805] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2805] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2805]] = 0;
              ip = 6242;
      end

       6242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 6] = localMem[2805];
              updateArrayLength(1, localMem[2798], 6);
              ip = 6243;
      end

       6243 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2806] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2806] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2806]] = 0;
              ip = 6244;
      end

       6244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 6] = localMem[2806];
              updateArrayLength(1, localMem[2801], 6);
              ip = 6245;
      end

       6245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2807] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6246;
      end

       6246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2808] = heapMem[localMem[2798]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6247;
      end

       6247 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2808] + 0 + i] = heapMem[NArea * localMem[2807] + 0 + i];
                  updateArrayLength(1, localMem[2808], 0 + i);
                end
              end
              ip = 6248;
      end

       6248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2809] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6249;
      end

       6249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2810] = heapMem[localMem[2798]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6250;
      end

       6250 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2810] + 0 + i] = heapMem[NArea * localMem[2809] + 0 + i];
                  updateArrayLength(1, localMem[2810], 0 + i);
                end
              end
              ip = 6251;
      end

       6251 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2811] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6252;
      end

       6252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2812] = heapMem[localMem[2798]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6253;
      end

       6253 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2813] = localMem[2748] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6254;
      end

       6254 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2813]) begin
                  heapMem[NArea * localMem[2812] + 0 + i] = heapMem[NArea * localMem[2811] + 0 + i];
                  updateArrayLength(1, localMem[2812], 0 + i);
                end
              end
              ip = 6255;
      end

       6255 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2814] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6256;
      end

       6256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2815] = heapMem[localMem[2801]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6257;
      end

       6257 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2815] + 0 + i] = heapMem[NArea * localMem[2814] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2815], 0 + i);
                end
              end
              ip = 6258;
      end

       6258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2816] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6259;
      end

       6259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2817] = heapMem[localMem[2801]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6260;
      end

       6260 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2817] + 0 + i] = heapMem[NArea * localMem[2816] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2817], 0 + i);
                end
              end
              ip = 6261;
      end

       6261 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2818] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6262;
      end

       6262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2819] = heapMem[localMem[2801]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6263;
      end

       6263 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2820] = localMem[2748] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6264;
      end

       6264 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2820]) begin
                  heapMem[NArea * localMem[2819] + 0 + i] = heapMem[NArea * localMem[2818] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2819], 0 + i);
                end
              end
              ip = 6265;
      end

       6265 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2821] = heapMem[localMem[2798]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6266;
      end

       6266 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2822] = localMem[2821] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6267;
      end

       6267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2823] = heapMem[localMem[2798]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6268;
      end

       6268 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6269;
      end

       6269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2824] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6270;
      end

       6270 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6271;
      end

       6271 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2824] >= localMem[2822] ? 6277 : 6272;
      end

       6272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2825] = heapMem[localMem[2823]*6 + localMem[2824]];
              updateArrayLength(2, 0, 0);
              ip = 6273;
      end

       6273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2825]*6 + 2] = localMem[2798];
              updateArrayLength(1, localMem[2825], 2);
              ip = 6274;
      end

       6274 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6275;
      end

       6275 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2824] = localMem[2824] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6276;
      end

       6276 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6270;
      end

       6277 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6278;
      end

       6278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2826] = heapMem[localMem[2801]*6 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6279;
      end

       6279 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2827] = localMem[2826] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6280;
      end

       6280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2828] = heapMem[localMem[2801]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6281;
      end

       6281 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6282;
      end

       6282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2829] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6283;
      end

       6283 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6284;
      end

       6284 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2829] >= localMem[2827] ? 6290 : 6285;
      end

       6285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2830] = heapMem[localMem[2828]*6 + localMem[2829]];
              updateArrayLength(2, 0, 0);
              ip = 6286;
      end

       6286 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2830]*6 + 2] = localMem[2801];
              updateArrayLength(1, localMem[2830], 2);
              ip = 6287;
      end

       6287 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6288;
      end

       6288 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2829] = localMem[2829] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6289;
      end

       6289 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6283;
      end

       6290 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6291;
      end

       6291 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6307;
      end

       6292 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6293;
      end

       6293 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2831] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2831] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2831]] = 0;
              ip = 6294;
      end

       6294 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2735]*6 + 6] = localMem[2831];
              updateArrayLength(1, localMem[2735], 6);
              ip = 6295;
      end

       6295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2832] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6296;
      end

       6296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2833] = heapMem[localMem[2798]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6297;
      end

       6297 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2833] + 0 + i] = heapMem[NArea * localMem[2832] + 0 + i];
                  updateArrayLength(1, localMem[2833], 0 + i);
                end
              end
              ip = 6298;
      end

       6298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2834] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6299;
      end

       6299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2835] = heapMem[localMem[2798]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6300;
      end

       6300 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2835] + 0 + i] = heapMem[NArea * localMem[2834] + 0 + i];
                  updateArrayLength(1, localMem[2835], 0 + i);
                end
              end
              ip = 6301;
      end

       6301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2836] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6302;
      end

       6302 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2837] = heapMem[localMem[2801]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6303;
      end

       6303 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2837] + 0 + i] = heapMem[NArea * localMem[2836] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2837], 0 + i);
                end
              end
              ip = 6304;
      end

       6304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2838] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6305;
      end

       6305 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2839] = heapMem[localMem[2801]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6306;
      end

       6306 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2748]) begin
                  heapMem[NArea * localMem[2839] + 0 + i] = heapMem[NArea * localMem[2838] + localMem[2749] + i];
                  updateArrayLength(1, localMem[2839], 0 + i);
                end
              end
              ip = 6307;
      end

       6307 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6308;
      end

       6308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2798]*6 + 2] = localMem[2735];
              updateArrayLength(1, localMem[2798], 2);
              ip = 6309;
      end

       6309 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2801]*6 + 2] = localMem[2735];
              updateArrayLength(1, localMem[2801], 2);
              ip = 6310;
      end

       6310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2840] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6311;
      end

       6311 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2841] = heapMem[localMem[2840]*6 + localMem[2748]];
              updateArrayLength(2, 0, 0);
              ip = 6312;
      end

       6312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2842] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6313;
      end

       6313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2843] = heapMem[localMem[2842]*6 + localMem[2748]];
              updateArrayLength(2, 0, 0);
              ip = 6314;
      end

       6314 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2844] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6315;
      end

       6315 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2844]*6 + 0] = localMem[2841];
              updateArrayLength(1, localMem[2844], 0);
              ip = 6316;
      end

       6316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2845] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6317;
      end

       6317 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2845]*6 + 0] = localMem[2843];
              updateArrayLength(1, localMem[2845], 0);
              ip = 6318;
      end

       6318 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2846] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6319;
      end

       6319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2846]*6 + 0] = localMem[2798];
              updateArrayLength(1, localMem[2846], 0);
              ip = 6320;
      end

       6320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2847] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6321;
      end

       6321 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2847]*6 + 1] = localMem[2801];
              updateArrayLength(1, localMem[2847], 1);
              ip = 6322;
      end

       6322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2735]*6 + 0] = 1;
              updateArrayLength(1, localMem[2735], 0);
              ip = 6323;
      end

       6323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2848] = heapMem[localMem[2735]*6 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6324;
      end

       6324 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2848]] = 1;
              ip = 6325;
      end

       6325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2849] = heapMem[localMem[2735]*6 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6326;
      end

       6326 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2849]] = 1;
              ip = 6327;
      end

       6327 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2850] = heapMem[localMem[2735]*6 + 6];
              updateArrayLength(2, 0, 0);
              ip = 6328;
      end

       6328 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2850]] = 2;
              ip = 6329;
      end

       6329 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6331;
      end

       6330 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6336;
      end

       6331 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6332;
      end

       6332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2744] = 1;
              updateArrayLength(2, 0, 0);
              ip = 6333;
      end

       6333 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6336;
      end

       6334 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6335;
      end

       6335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2744] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6336;
      end

       6336 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6337;
      end

       6337 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6338;
      end

       6338 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6339;
      end

       6339 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6340;
      end

       6340 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[2376]] = 0;
              freedArrays[freedArraysTop] = localMem[2376];
              freedArraysTop = freedArraysTop + 1;
              ip = 6341;
      end
      default: begin
        success  = 1;
        finished = 1;
      end
    endcase
    if (steps <=    492) clock <= ~ clock;                                      // Must be non sequential to fire the next iteration
    if (0) begin
      for(i = 0; i < 200; ++i) $write("%2d",   localMem[i]); $display("");
      for(i = 0; i < 200; ++i) $write("%2d",    heapMem[i]); $display("");
      for(i = 0; i < 200; ++i) $write("%2d", arraySizes[i]); $display("");
    end
  end
endmodule
