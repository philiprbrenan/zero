  parameter integer NInstructions = 1141;

  task startTest();                                                             // BTree: load code
    begin

      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;                                                                          // array
      code[   1] = 'h0000002000000000000000000000010000000000000120000000000000000000;                                                                          // label
      code[   2] = 'h0000001600000000000000000001210000000000000000000000000000000000;                                                                          // inSize
      code[   3] = 'h0000001800000000000004710003210000000000000121000000000000000000;                                                                          // jFalse
      code[   4] = 'h0000001500000000000000000002210000000000000000000000000000000000;                                                                          // in
      code[   5] = 'h0000001d00000000000000070004210000000000000221000000000000002000;                                                                          // jNe
      code[   6] = 'h0000000100000000000000000003210000000000000420000000000000000000;                                                                          // array
      code[   7] = 'h0000002300000000000000030002150000000000000320000000000000000000;                                                                          // mov
      code[   8] = 'h0000002300000000000000030003150000000000000020000000000000000000;                                                                          // mov
      code[   9] = 'h0000002300000000000000030000150000000000000020000000000000000000;                                                                          // mov
      code[  10] = 'h0000002300000000000000030001150000000000000020000000000000000000;                                                                          // mov
      code[  11] = 'h0000001f00000000000004670002210000000000000000000000000000000000;                                                                          // jmp
      code[  12] = 'h0000002000000000000000000000010000000000000420000000000000000000;                                                                          // label
      code[  13] = 'h0000001d000000000000041d0005210000000000000221000000000000012000;                                                                          // jNe
      code[  14] = 'h0000001500000000000000000004210000000000000000000000000000000000;                                                                          // in
      code[  15] = 'h0000001500000000000000000005210000000000000000000000000000000000;                                                                          // in
      code[  16] = 'h0000000100000000000000000006210000000000000320000000000000000000;                                                                          // array
      code[  17] = 'h0000002000000000000000000000010000000000000620000000000000000000;                                                                          // label
      code[  18] = 'h0000002300000000000000000007210000000003000315000000000000000000;                                                                          // mov
      code[  19] = 'h0000001d0000000000000013000a210000000000000721000000000000002000;                                                                          // jNe
      code[  20] = 'h0000000100000000000000000008210000000000000520000000000000000000;                                                                          // array
      code[  21] = 'h0000002300000000000000080000150000000000000120000000000000000000;                                                                          // mov
      code[  22] = 'h0000002300000000000000080002150000000000000020000000000000000000;                                                                          // mov
      code[  23] = 'h0000000100000000000000000009210000000000000620000000000000000000;                                                                          // array
      code[  24] = 'h0000002300000000000000080004150000000000000921000000000000000000;                                                                          // mov
      code[  25] = 'h000000010000000000000000000a210000000000000720000000000000000000;                                                                          // array
      code[  26] = 'h0000002300000000000000080005150000000000000a21000000000000000000;                                                                          // mov
      code[  27] = 'h0000002300000000000000080006150000000000000020000000000000000000;                                                                          // mov
      code[  28] = 'h0000002300000000000000080003150000000000000321000000000000000000;                                                                          // mov
      code[  29] = 'h0000000000000000000000030001150000000003000115000000000000012000;                                                                          // add
      code[  30] = 'h0000002300000000000000080001150000000003000115000000000000000000;                                                                          // mov
      code[  31] = 'h000000230000000000000000000b210000000008000415000000000000000000;                                                                          // mov
      code[  32] = 'h00000023000000000000000b0000150000000000000421000000000000000000;                                                                          // mov
      code[  33] = 'h000000230000000000000000000c210000000008000515000000000000000000;                                                                          // mov
      code[  34] = 'h00000023000000000000000c0000150000000000000521000000000000000000;                                                                          // mov
      code[  35] = 'h0000000000000000000000030000150000000003000015000000000000012000;                                                                          // add
      code[  36] = 'h0000002300000000000000030003150000000000000821000000000000000000;                                                                          // mov
      code[  37] = 'h0000001f00000000000004020009210000000000000000000000000000000000;                                                                          // jmp
      code[  38] = 'h0000002000000000000000000000010000000000000a20000000000000000000;                                                                          // label
      code[  39] = 'h000000230000000000000000000d210000000007000015000000000000000000;                                                                          // mov
      code[  40] = 'h000000230000000000000000000e210000000003000215000000000000000000;                                                                          // mov
      code[  41] = 'h000000190000000000000021000b210000000000000d210000000000000e2100;                                                                          // jGe
      code[  42] = 'h000000230000000000000000000f210000000007000215000000000000000000;                                                                          // mov
      code[  43] = 'h0000001d000000000000001e000c210000000000000f21000000000000002000;                                                                          // jNe
      code[  44] = 'h0000002600000000000000000010210000000007000615000000000000000000;                                                                          // not
      code[  45] = 'h00000017000000000000001b000d210000000000001021000000000000002000;                                                                          // jEq
      code[  46] = 'h0000002300000000000000000011210000000007000415000000000000000000;                                                                          // mov
      code[  47] = 'h0000000500000000000000000012210000000000001121000000000000042100;                                                                          // arrayIndex
      code[  48] = 'h000000170000000000000005000e210000000000001221000000000000002000;                                                                          // jEq
      code[  49] = 'h0000003900000000000000000012210000000000001221000000000000012000;                                                                          // subtract
      code[  50] = 'h0000002300000000000000000013210000000007000515000000000000000000;                                                                          // mov
      code[  51] = 'h0000002300000000000000130012160000000000000521000000000000000000;                                                                          // mov
      code[  52] = 'h0000001f00000000000003f30009210000000000000000000000000000000000;                                                                          // jmp
      code[  53] = 'h0000002000000000000000000000010000000000000e20000000000000000000;                                                                          // label
      code[  54] = 'h0000000200000000000000000014210000000000001121000000000000042100;                                                                          // arrayCountGreater
      code[  55] = 'h0000001d0000000000000008000f210000000000001421000000000000002000;                                                                          // jNe
      code[  56] = 'h0000002300000000000000000015210000000007000415000000000000000000;                                                                          // mov
      code[  57] = 'h000000230000000000000015000d160000000000000421000000000000000000;                                                                          // mov
      code[  58] = 'h0000002300000000000000000016210000000007000515000000000000000000;                                                                          // mov
      code[  59] = 'h000000230000000000000016000d160000000000000521000000000000000000;                                                                          // mov
      code[  60] = 'h0000000000000000000000070000150000000000000d21000000000000012000;                                                                          // add
      code[  61] = 'h0000000000000000000000030000150000000003000015000000000000012000;                                                                          // add
      code[  62] = 'h0000001f00000000000003e90009210000000000000000000000000000000000;                                                                          // jmp
      code[  63] = 'h0000002000000000000000000000010000000000000f20000000000000000000;                                                                          // label
      code[  64] = 'h0000000300000000000000000017210000000000001121000000000000042100;                                                                          // arrayCountLess
      code[  65] = 'h0000002300000000000000000018210000000007000415000000000000000000;                                                                          // mov
      code[  66] = 'h0000003800000000000000180017160000000000000421000000000000000000;                                                                          // shiftUp
      code[  67] = 'h0000002300000000000000000019210000000007000515000000000000000000;                                                                          // mov
      code[  68] = 'h0000003800000000000000190017160000000000000521000000000000000000;                                                                          // shiftUp
      code[  69] = 'h0000000000000000000000070000150000000007000015000000000000012000;                                                                          // add
      code[  70] = 'h0000000000000000000000030000150000000003000015000000000000012000;                                                                          // add
      code[  71] = 'h0000001f00000000000003e00009210000000000000000000000000000000000;                                                                          // jmp
      code[  72] = 'h0000002000000000000000000000010000000000000d20000000000000000000;                                                                          // label
      code[  73] = 'h0000002000000000000000000000010000000000000c20000000000000000000;                                                                          // label
      code[  74] = 'h0000002000000000000000000000010000000000000b20000000000000000000;                                                                          // label
      code[  75] = 'h000000230000000000000000001a210000000003000315000000000000000000;                                                                          // mov
      code[  76] = 'h0000002000000000000000000000010000000000001020000000000000000000;                                                                          // label
      code[  77] = 'h000000230000000000000000001c21000000001a000015000000000000000000;                                                                          // mov
      code[  78] = 'h000000230000000000000000001d21000000001a000315000000000000000000;                                                                          // mov
      code[  79] = 'h000000230000000000000000001e21000000001d000215000000000000000000;                                                                          // mov
      code[  80] = 'h0000001c00000000000000dc0012210000000000001c210000000000001e2100;                                                                          // jLt
      code[  81] = 'h000000230000000000000000001f210000000000001e21000000000000000000;                                                                          // mov
      code[  82] = 'h000000370000000000000000001f210000000000000120000000000000000000;                                                                          // shiftRight
      code[  83] = 'h0000000000000000000000000020210000000000001f21000000000000012000;                                                                          // add
      code[  84] = 'h000000230000000000000000002121000000001a000215000000000000000000;                                                                          // mov
      code[  85] = 'h0000001700000000000000610014210000000000002121000000000000002000;                                                                          // jEq
      code[  86] = 'h0000000100000000000000000022210000000000000520000000000000000000;                                                                          // array
      code[  87] = 'h0000002300000000000000220000150000000000001f21000000000000000000;                                                                          // mov
      code[  88] = 'h0000002300000000000000220002150000000000000020000000000000000000;                                                                          // mov
      code[  89] = 'h0000000100000000000000000023210000000000000620000000000000000000;                                                                          // array
      code[  90] = 'h0000002300000000000000220004150000000000002321000000000000000000;                                                                          // mov
      code[  91] = 'h0000000100000000000000000024210000000000000720000000000000000000;                                                                          // array
      code[  92] = 'h0000002300000000000000220005150000000000002421000000000000000000;                                                                          // mov
      code[  93] = 'h0000002300000000000000220006150000000000000020000000000000000000;                                                                          // mov
      code[  94] = 'h0000002300000000000000220003150000000000001d21000000000000000000;                                                                          // mov
      code[  95] = 'h00000000000000000000001d000115000000001d000115000000000000012000;                                                                          // add
      code[  96] = 'h000000230000000000000022000115000000001d000115000000000000000000;                                                                          // mov
      code[  97] = 'h000000260000000000000000002521000000001a000615000000000000000000;                                                                          // not
      code[  98] = 'h0000001d000000000000001d0015210000000000002521000000000000002000;                                                                          // jNe
      code[  99] = 'h0000000100000000000000000026210000000000000820000000000000000000;                                                                          // array
      code[ 100] = 'h0000002300000000000000220006150000000000002621000000000000000000;                                                                          // mov
      code[ 101] = 'h000000230000000000000000002721000000001a000415000000000000000000;                                                                          // mov
      code[ 102] = 'h0000002300000000000000000028210000000022000415000000000000000000;                                                                          // mov
      code[ 103] = 'h00000024000000000000002800001500000000270020160000000000001f2100;                                                                          // moveLong
      code[ 104] = 'h000000230000000000000000002921000000001a000515000000000000000000;                                                                          // mov
      code[ 105] = 'h000000230000000000000000002a210000000022000515000000000000000000;                                                                          // mov
      code[ 106] = 'h00000024000000000000002a00001500000000290020160000000000001f2100;                                                                          // moveLong
      code[ 107] = 'h000000230000000000000000002b21000000001a000615000000000000000000;                                                                          // mov
      code[ 108] = 'h000000230000000000000000002c210000000022000615000000000000000000;                                                                          // mov
      code[ 109] = 'h000000000000000000000000002d210000000000001f21000000000000012000;                                                                          // add
      code[ 110] = 'h00000024000000000000002c000015000000002b0020160000000000002d2100;                                                                          // moveLong
      code[ 111] = 'h000000230000000000000000002e210000000022000015000000000000000000;                                                                          // mov
      code[ 112] = 'h000000000000000000000000002f210000000000002e21000000000000012000;                                                                          // add
      code[ 113] = 'h0000002300000000000000000030210000000022000615000000000000000000;                                                                          // mov
      code[ 114] = 'h0000002000000000000000000000010000000000001720000000000000000000;                                                                          // label
      code[ 115] = 'h0000002300000000000000000031210000000000000020000000000000000000;                                                                          // mov
      code[ 116] = 'h0000002000000000000000000000010000000000001820000000000000000000;                                                                          // label
      code[ 117] = 'h000000190000000000000006001a2100000000000031210000000000002f2100;                                                                          // jGe
      code[ 118] = 'h0000002300000000000000000032210000000030003116000000000000000000;                                                                          // mov
      code[ 119] = 'h0000002300000000000000320002150000000000002221000000000000000000;                                                                          // mov
      code[ 120] = 'h0000002000000000000000000000010000000000001920000000000000000000;                                                                          // label
      code[ 121] = 'h0000000000000000000000000031210000000000003121000000000000012000;                                                                          // add
      code[ 122] = 'h0000001f00000000fffffffa0018210000000000000000000000000000000000;                                                                          // jmp
      code[ 123] = 'h0000002000000000000000000000010000000000001a20000000000000000000;                                                                          // label
      code[ 124] = 'h000000230000000000000000003321000000001a000615000000000000000000;                                                                          // mov
      code[ 125] = 'h0000003100000000000000000033210000000000002021000000000000082000;                                                                          // resize
      code[ 126] = 'h0000001f00000000000000080016210000000000000000000000000000000000;                                                                          // jmp
      code[ 127] = 'h0000002000000000000000000000010000000000001520000000000000000000;                                                                          // label
      code[ 128] = 'h000000230000000000000000003421000000001a000415000000000000000000;                                                                          // mov
      code[ 129] = 'h0000002300000000000000000035210000000022000415000000000000000000;                                                                          // mov
      code[ 130] = 'h00000024000000000000003500001500000000340020160000000000001f2100;                                                                          // moveLong
      code[ 131] = 'h000000230000000000000000003621000000001a000515000000000000000000;                                                                          // mov
      code[ 132] = 'h0000002300000000000000000037210000000022000515000000000000000000;                                                                          // mov
      code[ 133] = 'h00000024000000000000003700001500000000360020160000000000001f2100;                                                                          // moveLong
      code[ 134] = 'h0000002000000000000000000000010000000000001620000000000000000000;                                                                          // label
      code[ 135] = 'h00000023000000000000001a0000150000000000001f21000000000000000000;                                                                          // mov
      code[ 136] = 'h0000002300000000000000220002150000000000002121000000000000000000;                                                                          // mov
      code[ 137] = 'h0000002300000000000000000038210000000021000015000000000000000000;                                                                          // mov
      code[ 138] = 'h0000002300000000000000000039210000000021000615000000000000000000;                                                                          // mov
      code[ 139] = 'h000000230000000000000000003a210000000039003816000000000000000000;                                                                          // mov
      code[ 140] = 'h0000001d0000000000000013001b210000000000003a210000000000001a2100;                                                                          // jNe
      code[ 141] = 'h000000230000000000000000003b21000000001a000415000000000000000000;                                                                          // mov
      code[ 142] = 'h000000230000000000000000003c21000000003b001f16000000000000000000;                                                                          // mov
      code[ 143] = 'h000000230000000000000000003d210000000021000415000000000000000000;                                                                          // mov
      code[ 144] = 'h00000023000000000000003d0038160000000000003c21000000000000000000;                                                                          // mov
      code[ 145] = 'h000000230000000000000000003e21000000001a000515000000000000000000;                                                                          // mov
      code[ 146] = 'h000000230000000000000000003f21000000003e001f16000000000000000000;                                                                          // mov
      code[ 147] = 'h0000002300000000000000000040210000000021000515000000000000000000;                                                                          // mov
      code[ 148] = 'h0000002300000000000000400038160000000000003f21000000000000000000;                                                                          // mov
      code[ 149] = 'h000000230000000000000000004121000000001a000415000000000000000000;                                                                          // mov
      code[ 150] = 'h0000003100000000000000000041210000000000001f21000000000000062000;                                                                          // resize
      code[ 151] = 'h000000230000000000000000004221000000001a000515000000000000000000;                                                                          // mov
      code[ 152] = 'h0000003100000000000000000042210000000000001f21000000000000072000;                                                                          // resize
      code[ 153] = 'h0000000000000000000000000043210000000000003821000000000000012000;                                                                          // add
      code[ 154] = 'h0000002300000000000000210000150000000000004321000000000000000000;                                                                          // mov
      code[ 155] = 'h0000002300000000000000000044210000000021000615000000000000000000;                                                                          // mov
      code[ 156] = 'h0000002300000000000000440043160000000000002221000000000000000000;                                                                          // mov
      code[ 157] = 'h0000001f000000000000008c0011210000000000000000000000000000000000;                                                                          // jmp
      code[ 158] = 'h0000001f0000000000000017001c210000000000000000000000000000000000;                                                                          // jmp
      code[ 159] = 'h0000002000000000000000000000010000000000001b20000000000000000000;                                                                          // label
      code[ 160] = 'h0000000f00000000000000000000010000000000002121000000000000002000;                                                                          // assertNe
      code[ 161] = 'h0000002300000000000000000045210000000021000615000000000000000000;                                                                          // mov
      code[ 162] = 'h00000005000000000000000000462100000000000045210000000000001a2100;                                                                          // arrayIndex
      code[ 163] = 'h0000003900000000000000000046210000000000004621000000000000012000;                                                                          // subtract
      code[ 164] = 'h000000230000000000000000004721000000001a000415000000000000000000;                                                                          // mov
      code[ 165] = 'h0000002300000000000000000048210000000047001f16000000000000000000;                                                                          // mov
      code[ 166] = 'h000000230000000000000000004921000000001a000515000000000000000000;                                                                          // mov
      code[ 167] = 'h000000230000000000000000004a210000000049001f16000000000000000000;                                                                          // mov
      code[ 168] = 'h000000230000000000000000004b21000000001a000415000000000000000000;                                                                          // mov
      code[ 169] = 'h000000310000000000000000004b210000000000001f21000000000000062000;                                                                          // resize
      code[ 170] = 'h000000230000000000000000004c21000000001a000515000000000000000000;                                                                          // mov
      code[ 171] = 'h000000310000000000000000004c210000000000001f21000000000000072000;                                                                          // resize
      code[ 172] = 'h000000230000000000000000004d210000000021000415000000000000000000;                                                                          // mov
      code[ 173] = 'h00000038000000000000004d0046160000000000004821000000000000000000;                                                                          // shiftUp
      code[ 174] = 'h000000230000000000000000004e210000000021000515000000000000000000;                                                                          // mov
      code[ 175] = 'h00000038000000000000004e0046160000000000004a21000000000000000000;                                                                          // shiftUp
      code[ 176] = 'h000000230000000000000000004f210000000021000615000000000000000000;                                                                          // mov
      code[ 177] = 'h0000000000000000000000000050210000000000004621000000000000012000;                                                                          // add
      code[ 178] = 'h00000038000000000000004f0050160000000000002221000000000000000000;                                                                          // shiftUp
      code[ 179] = 'h0000000000000000000000210000150000000021000015000000000000012000;                                                                          // add
      code[ 180] = 'h0000001f00000000000000750011210000000000000000000000000000000000;                                                                          // jmp
      code[ 181] = 'h0000002000000000000000000000010000000000001c20000000000000000000;                                                                          // label
      code[ 182] = 'h0000002000000000000000000000010000000000001420000000000000000000;                                                                          // label
      code[ 183] = 'h0000000100000000000000000051210000000000000520000000000000000000;                                                                          // array
      code[ 184] = 'h0000002300000000000000510000150000000000001f21000000000000000000;                                                                          // mov
      code[ 185] = 'h0000002300000000000000510002150000000000000020000000000000000000;                                                                          // mov
      code[ 186] = 'h0000000100000000000000000052210000000000000620000000000000000000;                                                                          // array
      code[ 187] = 'h0000002300000000000000510004150000000000005221000000000000000000;                                                                          // mov
      code[ 188] = 'h0000000100000000000000000053210000000000000720000000000000000000;                                                                          // array
      code[ 189] = 'h0000002300000000000000510005150000000000005321000000000000000000;                                                                          // mov
      code[ 190] = 'h0000002300000000000000510006150000000000000020000000000000000000;                                                                          // mov
      code[ 191] = 'h0000002300000000000000510003150000000000001d21000000000000000000;                                                                          // mov
      code[ 192] = 'h00000000000000000000001d000115000000001d000115000000000000012000;                                                                          // add
      code[ 193] = 'h000000230000000000000051000115000000001d000115000000000000000000;                                                                          // mov
      code[ 194] = 'h0000000100000000000000000054210000000000000520000000000000000000;                                                                          // array
      code[ 195] = 'h0000002300000000000000540000150000000000001f21000000000000000000;                                                                          // mov
      code[ 196] = 'h0000002300000000000000540002150000000000000020000000000000000000;                                                                          // mov
      code[ 197] = 'h0000000100000000000000000055210000000000000620000000000000000000;                                                                          // array
      code[ 198] = 'h0000002300000000000000540004150000000000005521000000000000000000;                                                                          // mov
      code[ 199] = 'h0000000100000000000000000056210000000000000720000000000000000000;                                                                          // array
      code[ 200] = 'h0000002300000000000000540005150000000000005621000000000000000000;                                                                          // mov
      code[ 201] = 'h0000002300000000000000540006150000000000000020000000000000000000;                                                                          // mov
      code[ 202] = 'h0000002300000000000000540003150000000000001d21000000000000000000;                                                                          // mov
      code[ 203] = 'h00000000000000000000001d000115000000001d000115000000000000012000;                                                                          // add
      code[ 204] = 'h000000230000000000000054000115000000001d000115000000000000000000;                                                                          // mov
      code[ 205] = 'h000000260000000000000000005721000000001a000615000000000000000000;                                                                          // not
      code[ 206] = 'h0000001d0000000000000034001d210000000000005721000000000000002000;                                                                          // jNe
      code[ 207] = 'h0000000100000000000000000058210000000000000820000000000000000000;                                                                          // array
      code[ 208] = 'h0000002300000000000000510006150000000000005821000000000000000000;                                                                          // mov
      code[ 209] = 'h0000000100000000000000000059210000000000000820000000000000000000;                                                                          // array
      code[ 210] = 'h0000002300000000000000540006150000000000005921000000000000000000;                                                                          // mov
      code[ 211] = 'h000000230000000000000000005a21000000001a000415000000000000000000;                                                                          // mov
      code[ 212] = 'h000000230000000000000000005b210000000051000415000000000000000000;                                                                          // mov
      code[ 213] = 'h00000024000000000000005b000015000000005a0000150000000000001f2100;                                                                          // moveLong
      code[ 214] = 'h000000230000000000000000005c21000000001a000515000000000000000000;                                                                          // mov
      code[ 215] = 'h000000230000000000000000005d210000000051000515000000000000000000;                                                                          // mov
      code[ 216] = 'h00000024000000000000005d000015000000005c0000150000000000001f2100;                                                                          // moveLong
      code[ 217] = 'h000000230000000000000000005e21000000001a000615000000000000000000;                                                                          // mov
      code[ 218] = 'h000000230000000000000000005f210000000051000615000000000000000000;                                                                          // mov
      code[ 219] = 'h0000000000000000000000000060210000000000001f21000000000000012000;                                                                          // add
      code[ 220] = 'h00000024000000000000005f000015000000005e000015000000000000602100;                                                                          // moveLong
      code[ 221] = 'h000000230000000000000000006121000000001a000415000000000000000000;                                                                          // mov
      code[ 222] = 'h0000002300000000000000000062210000000054000415000000000000000000;                                                                          // mov
      code[ 223] = 'h00000024000000000000006200001500000000610020160000000000001f2100;                                                                          // moveLong
      code[ 224] = 'h000000230000000000000000006321000000001a000515000000000000000000;                                                                          // mov
      code[ 225] = 'h0000002300000000000000000064210000000054000515000000000000000000;                                                                          // mov
      code[ 226] = 'h00000024000000000000006400001500000000630020160000000000001f2100;                                                                          // moveLong
      code[ 227] = 'h000000230000000000000000006521000000001a000615000000000000000000;                                                                          // mov
      code[ 228] = 'h0000002300000000000000000066210000000054000615000000000000000000;                                                                          // mov
      code[ 229] = 'h0000000000000000000000000067210000000000001f21000000000000012000;                                                                          // add
      code[ 230] = 'h0000002400000000000000660000150000000065002016000000000000672100;                                                                          // moveLong
      code[ 231] = 'h0000002300000000000000000068210000000051000015000000000000000000;                                                                          // mov
      code[ 232] = 'h0000000000000000000000000069210000000000006821000000000000012000;                                                                          // add
      code[ 233] = 'h000000230000000000000000006a210000000051000615000000000000000000;                                                                          // mov
      code[ 234] = 'h0000002000000000000000000000010000000000001f20000000000000000000;                                                                          // label
      code[ 235] = 'h000000230000000000000000006b210000000000000020000000000000000000;                                                                          // mov
      code[ 236] = 'h0000002000000000000000000000010000000000002020000000000000000000;                                                                          // label
      code[ 237] = 'h0000001900000000000000060022210000000000006b21000000000000692100;                                                                          // jGe
      code[ 238] = 'h000000230000000000000000006c21000000006a006b16000000000000000000;                                                                          // mov
      code[ 239] = 'h00000023000000000000006c0002150000000000005121000000000000000000;                                                                          // mov
      code[ 240] = 'h0000002000000000000000000000010000000000002120000000000000000000;                                                                          // label
      code[ 241] = 'h000000000000000000000000006b210000000000006b21000000000000012000;                                                                          // add
      code[ 242] = 'h0000001f00000000fffffffa0020210000000000000000000000000000000000;                                                                          // jmp
      code[ 243] = 'h0000002000000000000000000000010000000000002220000000000000000000;                                                                          // label
      code[ 244] = 'h000000230000000000000000006d210000000054000015000000000000000000;                                                                          // mov
      code[ 245] = 'h000000000000000000000000006e210000000000006d21000000000000012000;                                                                          // add
      code[ 246] = 'h000000230000000000000000006f210000000054000615000000000000000000;                                                                          // mov
      code[ 247] = 'h0000002000000000000000000000010000000000002320000000000000000000;                                                                          // label
      code[ 248] = 'h0000002300000000000000000070210000000000000020000000000000000000;                                                                          // mov
      code[ 249] = 'h0000002000000000000000000000010000000000002420000000000000000000;                                                                          // label
      code[ 250] = 'h00000019000000000000000600262100000000000070210000000000006e2100;                                                                          // jGe
      code[ 251] = 'h000000230000000000000000007121000000006f007016000000000000000000;                                                                          // mov
      code[ 252] = 'h0000002300000000000000710002150000000000005421000000000000000000;                                                                          // mov
      code[ 253] = 'h0000002000000000000000000000010000000000002520000000000000000000;                                                                          // label
      code[ 254] = 'h0000000000000000000000000070210000000000007021000000000000012000;                                                                          // add
      code[ 255] = 'h0000001f00000000fffffffa0024210000000000000000000000000000000000;                                                                          // jmp
      code[ 256] = 'h0000002000000000000000000000010000000000002620000000000000000000;                                                                          // label
      code[ 257] = 'h0000001f0000000000000010001e210000000000000000000000000000000000;                                                                          // jmp
      code[ 258] = 'h0000002000000000000000000000010000000000001d20000000000000000000;                                                                          // label
      code[ 259] = 'h0000000100000000000000000072210000000000000820000000000000000000;                                                                          // array
      code[ 260] = 'h00000023000000000000001a0006150000000000007221000000000000000000;                                                                          // mov
      code[ 261] = 'h000000230000000000000000007321000000001a000415000000000000000000;                                                                          // mov
      code[ 262] = 'h0000002300000000000000000074210000000051000415000000000000000000;                                                                          // mov
      code[ 263] = 'h00000024000000000000007400001500000000730000150000000000001f2100;                                                                          // moveLong
      code[ 264] = 'h000000230000000000000000007521000000001a000515000000000000000000;                                                                          // mov
      code[ 265] = 'h0000002300000000000000000076210000000051000515000000000000000000;                                                                          // mov
      code[ 266] = 'h00000024000000000000007600001500000000750000150000000000001f2100;                                                                          // moveLong
      code[ 267] = 'h000000230000000000000000007721000000001a000415000000000000000000;                                                                          // mov
      code[ 268] = 'h0000002300000000000000000078210000000054000415000000000000000000;                                                                          // mov
      code[ 269] = 'h00000024000000000000007800001500000000770020160000000000001f2100;                                                                          // moveLong
      code[ 270] = 'h000000230000000000000000007921000000001a000515000000000000000000;                                                                          // mov
      code[ 271] = 'h000000230000000000000000007a210000000054000515000000000000000000;                                                                          // mov
      code[ 272] = 'h00000024000000000000007a00001500000000790020160000000000001f2100;                                                                          // moveLong
      code[ 273] = 'h0000002000000000000000000000010000000000001e20000000000000000000;                                                                          // label
      code[ 274] = 'h0000002300000000000000510002150000000000001a21000000000000000000;                                                                          // mov
      code[ 275] = 'h0000002300000000000000540002150000000000001a21000000000000000000;                                                                          // mov
      code[ 276] = 'h000000230000000000000000007b21000000001a000415000000000000000000;                                                                          // mov
      code[ 277] = 'h000000230000000000000000007c21000000007b001f16000000000000000000;                                                                          // mov
      code[ 278] = 'h000000230000000000000000007d21000000001a000515000000000000000000;                                                                          // mov
      code[ 279] = 'h000000230000000000000000007e21000000007d001f16000000000000000000;                                                                          // mov
      code[ 280] = 'h000000230000000000000000007f21000000001a000415000000000000000000;                                                                          // mov
      code[ 281] = 'h00000023000000000000007f0000150000000000007c21000000000000000000;                                                                          // mov
      code[ 282] = 'h000000230000000000000000008021000000001a000515000000000000000000;                                                                          // mov
      code[ 283] = 'h0000002300000000000000800000150000000000007e21000000000000000000;                                                                          // mov
      code[ 284] = 'h000000230000000000000000008121000000001a000615000000000000000000;                                                                          // mov
      code[ 285] = 'h0000002300000000000000810000150000000000005121000000000000000000;                                                                          // mov
      code[ 286] = 'h000000230000000000000000008221000000001a000615000000000000000000;                                                                          // mov
      code[ 287] = 'h0000002300000000000000820001150000000000005421000000000000000000;                                                                          // mov
      code[ 288] = 'h00000023000000000000001a0000150000000000000120000000000000000000;                                                                          // mov
      code[ 289] = 'h000000230000000000000000008321000000001a000415000000000000000000;                                                                          // mov
      code[ 290] = 'h0000003100000000000000000083210000000000000120000000000000062000;                                                                          // resize
      code[ 291] = 'h000000230000000000000000008421000000001a000515000000000000000000;                                                                          // mov
      code[ 292] = 'h0000003100000000000000000084210000000000000120000000000000072000;                                                                          // resize
      code[ 293] = 'h000000230000000000000000008521000000001a000615000000000000000000;                                                                          // mov
      code[ 294] = 'h0000003100000000000000000085210000000000000220000000000000082000;                                                                          // resize
      code[ 295] = 'h0000001f00000000000000020011210000000000000000000000000000000000;                                                                          // jmp
      code[ 296] = 'h0000001f00000000000000060013210000000000000000000000000000000000;                                                                          // jmp
      code[ 297] = 'h0000002000000000000000000000010000000000001120000000000000000000;                                                                          // label
      code[ 298] = 'h000000230000000000000000001b210000000000000120000000000000000000;                                                                          // mov
      code[ 299] = 'h0000001f00000000000000030013210000000000000000000000000000000000;                                                                          // jmp
      code[ 300] = 'h0000002000000000000000000000010000000000001220000000000000000000;                                                                          // label
      code[ 301] = 'h000000230000000000000000001b210000000000000020000000000000000000;                                                                          // mov
      code[ 302] = 'h0000002000000000000000000000010000000000001320000000000000000000;                                                                          // label
      code[ 303] = 'h0000002000000000000000000000010000000000002720000000000000000000;                                                                          // label
      code[ 304] = 'h0000002000000000000000000000010000000000002b20000000000000000000;                                                                          // label
      code[ 305] = 'h0000002300000000000000000086210000000000000020000000000000000000;                                                                          // mov
      code[ 306] = 'h0000002000000000000000000000010000000000002c20000000000000000000;                                                                          // label
      code[ 307] = 'h0000001900000000000001f2002e210000000000008621000000000000632000;                                                                          // jGe
      code[ 308] = 'h000000230000000000000000008721000000001a000015000000000000000000;                                                                          // mov
      code[ 309] = 'h0000003900000000000000000088210000000000008721000000000000012000;                                                                          // subtract
      code[ 310] = 'h000000230000000000000000008921000000001a000415000000000000000000;                                                                          // mov
      code[ 311] = 'h000000230000000000000000008a210000000089008816000000000000000000;                                                                          // mov
      code[ 312] = 'h0000001b00000000000000f1002f2100000000000004210000000000008a2100;                                                                          // jLe
      code[ 313] = 'h000000260000000000000000008b21000000001a000615000000000000000000;                                                                          // not
      code[ 314] = 'h0000001700000000000000050030210000000000008b21000000000000002000;                                                                          // jEq
      code[ 315] = 'h0000002300000000000000060000150000000000001a21000000000000000000;                                                                          // mov
      code[ 316] = 'h0000002300000000000000060001150000000000000220000000000000000000;                                                                          // mov
      code[ 317] = 'h0000003900000000000000060002150000000000008721000000000000012000;                                                                          // subtract
      code[ 318] = 'h0000001f00000000000001eb002a210000000000000000000000000000000000;                                                                          // jmp
      code[ 319] = 'h0000002000000000000000000000010000000000003020000000000000000000;                                                                          // label
      code[ 320] = 'h000000230000000000000000008c21000000001a000615000000000000000000;                                                                          // mov
      code[ 321] = 'h000000230000000000000000008d21000000008c008716000000000000000000;                                                                          // mov
      code[ 322] = 'h0000002000000000000000000000010000000000003120000000000000000000;                                                                          // label
      code[ 323] = 'h000000230000000000000000008f21000000008d000015000000000000000000;                                                                          // mov
      code[ 324] = 'h000000230000000000000000009021000000008d000315000000000000000000;                                                                          // mov
      code[ 325] = 'h0000002300000000000000000091210000000090000215000000000000000000;                                                                          // mov
      code[ 326] = 'h0000001c00000000000000dc0033210000000000008f21000000000000912100;                                                                          // jLt
      code[ 327] = 'h0000002300000000000000000092210000000000009121000000000000000000;                                                                          // mov
      code[ 328] = 'h0000003700000000000000000092210000000000000120000000000000000000;                                                                          // shiftRight
      code[ 329] = 'h0000000000000000000000000093210000000000009221000000000000012000;                                                                          // add
      code[ 330] = 'h000000230000000000000000009421000000008d000215000000000000000000;                                                                          // mov
      code[ 331] = 'h0000001700000000000000610035210000000000009421000000000000002000;                                                                          // jEq
      code[ 332] = 'h0000000100000000000000000095210000000000000520000000000000000000;                                                                          // array
      code[ 333] = 'h0000002300000000000000950000150000000000009221000000000000000000;                                                                          // mov
      code[ 334] = 'h0000002300000000000000950002150000000000000020000000000000000000;                                                                          // mov
      code[ 335] = 'h0000000100000000000000000096210000000000000620000000000000000000;                                                                          // array
      code[ 336] = 'h0000002300000000000000950004150000000000009621000000000000000000;                                                                          // mov
      code[ 337] = 'h0000000100000000000000000097210000000000000720000000000000000000;                                                                          // array
      code[ 338] = 'h0000002300000000000000950005150000000000009721000000000000000000;                                                                          // mov
      code[ 339] = 'h0000002300000000000000950006150000000000000020000000000000000000;                                                                          // mov
      code[ 340] = 'h0000002300000000000000950003150000000000009021000000000000000000;                                                                          // mov
      code[ 341] = 'h0000000000000000000000900001150000000090000115000000000000012000;                                                                          // add
      code[ 342] = 'h0000002300000000000000950001150000000090000115000000000000000000;                                                                          // mov
      code[ 343] = 'h000000260000000000000000009821000000008d000615000000000000000000;                                                                          // not
      code[ 344] = 'h0000001d000000000000001d0036210000000000009821000000000000002000;                                                                          // jNe
      code[ 345] = 'h0000000100000000000000000099210000000000000820000000000000000000;                                                                          // array
      code[ 346] = 'h0000002300000000000000950006150000000000009921000000000000000000;                                                                          // mov
      code[ 347] = 'h000000230000000000000000009a21000000008d000415000000000000000000;                                                                          // mov
      code[ 348] = 'h000000230000000000000000009b210000000095000415000000000000000000;                                                                          // mov
      code[ 349] = 'h00000024000000000000009b000015000000009a009316000000000000922100;                                                                          // moveLong
      code[ 350] = 'h000000230000000000000000009c21000000008d000515000000000000000000;                                                                          // mov
      code[ 351] = 'h000000230000000000000000009d210000000095000515000000000000000000;                                                                          // mov
      code[ 352] = 'h00000024000000000000009d000015000000009c009316000000000000922100;                                                                          // moveLong
      code[ 353] = 'h000000230000000000000000009e21000000008d000615000000000000000000;                                                                          // mov
      code[ 354] = 'h000000230000000000000000009f210000000095000615000000000000000000;                                                                          // mov
      code[ 355] = 'h00000000000000000000000000a0210000000000009221000000000000012000;                                                                          // add
      code[ 356] = 'h00000024000000000000009f000015000000009e009316000000000000a02100;                                                                          // moveLong
      code[ 357] = 'h00000023000000000000000000a1210000000095000015000000000000000000;                                                                          // mov
      code[ 358] = 'h00000000000000000000000000a221000000000000a121000000000000012000;                                                                          // add
      code[ 359] = 'h00000023000000000000000000a3210000000095000615000000000000000000;                                                                          // mov
      code[ 360] = 'h0000002000000000000000000000010000000000003820000000000000000000;                                                                          // label
      code[ 361] = 'h00000023000000000000000000a4210000000000000020000000000000000000;                                                                          // mov
      code[ 362] = 'h0000002000000000000000000000010000000000003920000000000000000000;                                                                          // label
      code[ 363] = 'h000000190000000000000006003b21000000000000a421000000000000a22100;                                                                          // jGe
      code[ 364] = 'h00000023000000000000000000a52100000000a300a416000000000000000000;                                                                          // mov
      code[ 365] = 'h0000002300000000000000a50002150000000000009521000000000000000000;                                                                          // mov
      code[ 366] = 'h0000002000000000000000000000010000000000003a20000000000000000000;                                                                          // label
      code[ 367] = 'h00000000000000000000000000a421000000000000a421000000000000012000;                                                                          // add
      code[ 368] = 'h0000001f00000000fffffffa0039210000000000000000000000000000000000;                                                                          // jmp
      code[ 369] = 'h0000002000000000000000000000010000000000003b20000000000000000000;                                                                          // label
      code[ 370] = 'h00000023000000000000000000a621000000008d000615000000000000000000;                                                                          // mov
      code[ 371] = 'h00000031000000000000000000a6210000000000009321000000000000082000;                                                                          // resize
      code[ 372] = 'h0000001f00000000000000080037210000000000000000000000000000000000;                                                                          // jmp
      code[ 373] = 'h0000002000000000000000000000010000000000003620000000000000000000;                                                                          // label
      code[ 374] = 'h00000023000000000000000000a721000000008d000415000000000000000000;                                                                          // mov
      code[ 375] = 'h00000023000000000000000000a8210000000095000415000000000000000000;                                                                          // mov
      code[ 376] = 'h0000002400000000000000a800001500000000a7009316000000000000922100;                                                                          // moveLong
      code[ 377] = 'h00000023000000000000000000a921000000008d000515000000000000000000;                                                                          // mov
      code[ 378] = 'h00000023000000000000000000aa210000000095000515000000000000000000;                                                                          // mov
      code[ 379] = 'h0000002400000000000000aa00001500000000a9009316000000000000922100;                                                                          // moveLong
      code[ 380] = 'h0000002000000000000000000000010000000000003720000000000000000000;                                                                          // label
      code[ 381] = 'h00000023000000000000008d0000150000000000009221000000000000000000;                                                                          // mov
      code[ 382] = 'h0000002300000000000000950002150000000000009421000000000000000000;                                                                          // mov
      code[ 383] = 'h00000023000000000000000000ab210000000094000015000000000000000000;                                                                          // mov
      code[ 384] = 'h00000023000000000000000000ac210000000094000615000000000000000000;                                                                          // mov
      code[ 385] = 'h00000023000000000000000000ad2100000000ac00ab16000000000000000000;                                                                          // mov
      code[ 386] = 'h0000001d0000000000000013003c21000000000000ad210000000000008d2100;                                                                          // jNe
      code[ 387] = 'h00000023000000000000000000ae21000000008d000415000000000000000000;                                                                          // mov
      code[ 388] = 'h00000023000000000000000000af2100000000ae009216000000000000000000;                                                                          // mov
      code[ 389] = 'h00000023000000000000000000b0210000000094000415000000000000000000;                                                                          // mov
      code[ 390] = 'h0000002300000000000000b000ab16000000000000af21000000000000000000;                                                                          // mov
      code[ 391] = 'h00000023000000000000000000b121000000008d000515000000000000000000;                                                                          // mov
      code[ 392] = 'h00000023000000000000000000b22100000000b1009216000000000000000000;                                                                          // mov
      code[ 393] = 'h00000023000000000000000000b3210000000094000515000000000000000000;                                                                          // mov
      code[ 394] = 'h0000002300000000000000b300ab16000000000000b221000000000000000000;                                                                          // mov
      code[ 395] = 'h00000023000000000000000000b421000000008d000415000000000000000000;                                                                          // mov
      code[ 396] = 'h00000031000000000000000000b4210000000000009221000000000000062000;                                                                          // resize
      code[ 397] = 'h00000023000000000000000000b521000000008d000515000000000000000000;                                                                          // mov
      code[ 398] = 'h00000031000000000000000000b5210000000000009221000000000000072000;                                                                          // resize
      code[ 399] = 'h00000000000000000000000000b621000000000000ab21000000000000012000;                                                                          // add
      code[ 400] = 'h000000230000000000000094000015000000000000b621000000000000000000;                                                                          // mov
      code[ 401] = 'h00000023000000000000000000b7210000000094000615000000000000000000;                                                                          // mov
      code[ 402] = 'h0000002300000000000000b700b6160000000000009521000000000000000000;                                                                          // mov
      code[ 403] = 'h0000001f000000000000008c0032210000000000000000000000000000000000;                                                                          // jmp
      code[ 404] = 'h0000001f0000000000000017003d210000000000000000000000000000000000;                                                                          // jmp
      code[ 405] = 'h0000002000000000000000000000010000000000003c20000000000000000000;                                                                          // label
      code[ 406] = 'h0000000f00000000000000000000010000000000009421000000000000002000;                                                                          // assertNe
      code[ 407] = 'h00000023000000000000000000b8210000000094000615000000000000000000;                                                                          // mov
      code[ 408] = 'h00000005000000000000000000b921000000000000b8210000000000008d2100;                                                                          // arrayIndex
      code[ 409] = 'h00000039000000000000000000b921000000000000b921000000000000012000;                                                                          // subtract
      code[ 410] = 'h00000023000000000000000000ba21000000008d000415000000000000000000;                                                                          // mov
      code[ 411] = 'h00000023000000000000000000bb2100000000ba009216000000000000000000;                                                                          // mov
      code[ 412] = 'h00000023000000000000000000bc21000000008d000515000000000000000000;                                                                          // mov
      code[ 413] = 'h00000023000000000000000000bd2100000000bc009216000000000000000000;                                                                          // mov
      code[ 414] = 'h00000023000000000000000000be21000000008d000415000000000000000000;                                                                          // mov
      code[ 415] = 'h00000031000000000000000000be210000000000009221000000000000062000;                                                                          // resize
      code[ 416] = 'h00000023000000000000000000bf21000000008d000515000000000000000000;                                                                          // mov
      code[ 417] = 'h00000031000000000000000000bf210000000000009221000000000000072000;                                                                          // resize
      code[ 418] = 'h00000023000000000000000000c0210000000094000415000000000000000000;                                                                          // mov
      code[ 419] = 'h0000003800000000000000c000b916000000000000bb21000000000000000000;                                                                          // shiftUp
      code[ 420] = 'h00000023000000000000000000c1210000000094000515000000000000000000;                                                                          // mov
      code[ 421] = 'h0000003800000000000000c100b916000000000000bd21000000000000000000;                                                                          // shiftUp
      code[ 422] = 'h00000023000000000000000000c2210000000094000615000000000000000000;                                                                          // mov
      code[ 423] = 'h00000000000000000000000000c321000000000000b921000000000000012000;                                                                          // add
      code[ 424] = 'h0000003800000000000000c200c3160000000000009521000000000000000000;                                                                          // shiftUp
      code[ 425] = 'h0000000000000000000000940000150000000094000015000000000000012000;                                                                          // add
      code[ 426] = 'h0000001f00000000000000750032210000000000000000000000000000000000;                                                                          // jmp
      code[ 427] = 'h0000002000000000000000000000010000000000003d20000000000000000000;                                                                          // label
      code[ 428] = 'h0000002000000000000000000000010000000000003520000000000000000000;                                                                          // label
      code[ 429] = 'h00000001000000000000000000c4210000000000000520000000000000000000;                                                                          // array
      code[ 430] = 'h0000002300000000000000c40000150000000000009221000000000000000000;                                                                          // mov
      code[ 431] = 'h0000002300000000000000c40002150000000000000020000000000000000000;                                                                          // mov
      code[ 432] = 'h00000001000000000000000000c5210000000000000620000000000000000000;                                                                          // array
      code[ 433] = 'h0000002300000000000000c4000415000000000000c521000000000000000000;                                                                          // mov
      code[ 434] = 'h00000001000000000000000000c6210000000000000720000000000000000000;                                                                          // array
      code[ 435] = 'h0000002300000000000000c4000515000000000000c621000000000000000000;                                                                          // mov
      code[ 436] = 'h0000002300000000000000c40006150000000000000020000000000000000000;                                                                          // mov
      code[ 437] = 'h0000002300000000000000c40003150000000000009021000000000000000000;                                                                          // mov
      code[ 438] = 'h0000000000000000000000900001150000000090000115000000000000012000;                                                                          // add
      code[ 439] = 'h0000002300000000000000c40001150000000090000115000000000000000000;                                                                          // mov
      code[ 440] = 'h00000001000000000000000000c7210000000000000520000000000000000000;                                                                          // array
      code[ 441] = 'h0000002300000000000000c70000150000000000009221000000000000000000;                                                                          // mov
      code[ 442] = 'h0000002300000000000000c70002150000000000000020000000000000000000;                                                                          // mov
      code[ 443] = 'h00000001000000000000000000c8210000000000000620000000000000000000;                                                                          // array
      code[ 444] = 'h0000002300000000000000c7000415000000000000c821000000000000000000;                                                                          // mov
      code[ 445] = 'h00000001000000000000000000c9210000000000000720000000000000000000;                                                                          // array
      code[ 446] = 'h0000002300000000000000c7000515000000000000c921000000000000000000;                                                                          // mov
      code[ 447] = 'h0000002300000000000000c70006150000000000000020000000000000000000;                                                                          // mov
      code[ 448] = 'h0000002300000000000000c70003150000000000009021000000000000000000;                                                                          // mov
      code[ 449] = 'h0000000000000000000000900001150000000090000115000000000000012000;                                                                          // add
      code[ 450] = 'h0000002300000000000000c70001150000000090000115000000000000000000;                                                                          // mov
      code[ 451] = 'h00000026000000000000000000ca21000000008d000615000000000000000000;                                                                          // not
      code[ 452] = 'h0000001d0000000000000034003e21000000000000ca21000000000000002000;                                                                          // jNe
      code[ 453] = 'h00000001000000000000000000cb210000000000000820000000000000000000;                                                                          // array
      code[ 454] = 'h0000002300000000000000c4000615000000000000cb21000000000000000000;                                                                          // mov
      code[ 455] = 'h00000001000000000000000000cc210000000000000820000000000000000000;                                                                          // array
      code[ 456] = 'h0000002300000000000000c7000615000000000000cc21000000000000000000;                                                                          // mov
      code[ 457] = 'h00000023000000000000000000cd21000000008d000415000000000000000000;                                                                          // mov
      code[ 458] = 'h00000023000000000000000000ce2100000000c4000415000000000000000000;                                                                          // mov
      code[ 459] = 'h0000002400000000000000ce00001500000000cd000015000000000000922100;                                                                          // moveLong
      code[ 460] = 'h00000023000000000000000000cf21000000008d000515000000000000000000;                                                                          // mov
      code[ 461] = 'h00000023000000000000000000d02100000000c4000515000000000000000000;                                                                          // mov
      code[ 462] = 'h0000002400000000000000d000001500000000cf000015000000000000922100;                                                                          // moveLong
      code[ 463] = 'h00000023000000000000000000d121000000008d000615000000000000000000;                                                                          // mov
      code[ 464] = 'h00000023000000000000000000d22100000000c4000615000000000000000000;                                                                          // mov
      code[ 465] = 'h00000000000000000000000000d3210000000000009221000000000000012000;                                                                          // add
      code[ 466] = 'h0000002400000000000000d200001500000000d1000015000000000000d32100;                                                                          // moveLong
      code[ 467] = 'h00000023000000000000000000d421000000008d000415000000000000000000;                                                                          // mov
      code[ 468] = 'h00000023000000000000000000d52100000000c7000415000000000000000000;                                                                          // mov
      code[ 469] = 'h0000002400000000000000d500001500000000d4009316000000000000922100;                                                                          // moveLong
      code[ 470] = 'h00000023000000000000000000d621000000008d000515000000000000000000;                                                                          // mov
      code[ 471] = 'h00000023000000000000000000d72100000000c7000515000000000000000000;                                                                          // mov
      code[ 472] = 'h0000002400000000000000d700001500000000d6009316000000000000922100;                                                                          // moveLong
      code[ 473] = 'h00000023000000000000000000d821000000008d000615000000000000000000;                                                                          // mov
      code[ 474] = 'h00000023000000000000000000d92100000000c7000615000000000000000000;                                                                          // mov
      code[ 475] = 'h00000000000000000000000000da210000000000009221000000000000012000;                                                                          // add
      code[ 476] = 'h0000002400000000000000d900001500000000d8009316000000000000da2100;                                                                          // moveLong
      code[ 477] = 'h00000023000000000000000000db2100000000c4000015000000000000000000;                                                                          // mov
      code[ 478] = 'h00000000000000000000000000dc21000000000000db21000000000000012000;                                                                          // add
      code[ 479] = 'h00000023000000000000000000dd2100000000c4000615000000000000000000;                                                                          // mov
      code[ 480] = 'h0000002000000000000000000000010000000000004020000000000000000000;                                                                          // label
      code[ 481] = 'h00000023000000000000000000de210000000000000020000000000000000000;                                                                          // mov
      code[ 482] = 'h0000002000000000000000000000010000000000004120000000000000000000;                                                                          // label
      code[ 483] = 'h000000190000000000000006004321000000000000de21000000000000dc2100;                                                                          // jGe
      code[ 484] = 'h00000023000000000000000000df2100000000dd00de16000000000000000000;                                                                          // mov
      code[ 485] = 'h0000002300000000000000df000215000000000000c421000000000000000000;                                                                          // mov
      code[ 486] = 'h0000002000000000000000000000010000000000004220000000000000000000;                                                                          // label
      code[ 487] = 'h00000000000000000000000000de21000000000000de21000000000000012000;                                                                          // add
      code[ 488] = 'h0000001f00000000fffffffa0041210000000000000000000000000000000000;                                                                          // jmp
      code[ 489] = 'h0000002000000000000000000000010000000000004320000000000000000000;                                                                          // label
      code[ 490] = 'h00000023000000000000000000e02100000000c7000015000000000000000000;                                                                          // mov
      code[ 491] = 'h00000000000000000000000000e121000000000000e021000000000000012000;                                                                          // add
      code[ 492] = 'h00000023000000000000000000e22100000000c7000615000000000000000000;                                                                          // mov
      code[ 493] = 'h0000002000000000000000000000010000000000004420000000000000000000;                                                                          // label
      code[ 494] = 'h00000023000000000000000000e3210000000000000020000000000000000000;                                                                          // mov
      code[ 495] = 'h0000002000000000000000000000010000000000004520000000000000000000;                                                                          // label
      code[ 496] = 'h000000190000000000000006004721000000000000e321000000000000e12100;                                                                          // jGe
      code[ 497] = 'h00000023000000000000000000e42100000000e200e316000000000000000000;                                                                          // mov
      code[ 498] = 'h0000002300000000000000e4000215000000000000c721000000000000000000;                                                                          // mov
      code[ 499] = 'h0000002000000000000000000000010000000000004620000000000000000000;                                                                          // label
      code[ 500] = 'h00000000000000000000000000e321000000000000e321000000000000012000;                                                                          // add
      code[ 501] = 'h0000001f00000000fffffffa0045210000000000000000000000000000000000;                                                                          // jmp
      code[ 502] = 'h0000002000000000000000000000010000000000004720000000000000000000;                                                                          // label
      code[ 503] = 'h0000001f0000000000000010003f210000000000000000000000000000000000;                                                                          // jmp
      code[ 504] = 'h0000002000000000000000000000010000000000003e20000000000000000000;                                                                          // label
      code[ 505] = 'h00000001000000000000000000e5210000000000000820000000000000000000;                                                                          // array
      code[ 506] = 'h00000023000000000000008d000615000000000000e521000000000000000000;                                                                          // mov
      code[ 507] = 'h00000023000000000000000000e621000000008d000415000000000000000000;                                                                          // mov
      code[ 508] = 'h00000023000000000000000000e72100000000c4000415000000000000000000;                                                                          // mov
      code[ 509] = 'h0000002400000000000000e700001500000000e6000015000000000000922100;                                                                          // moveLong
      code[ 510] = 'h00000023000000000000000000e821000000008d000515000000000000000000;                                                                          // mov
      code[ 511] = 'h00000023000000000000000000e92100000000c4000515000000000000000000;                                                                          // mov
      code[ 512] = 'h0000002400000000000000e900001500000000e8000015000000000000922100;                                                                          // moveLong
      code[ 513] = 'h00000023000000000000000000ea21000000008d000415000000000000000000;                                                                          // mov
      code[ 514] = 'h00000023000000000000000000eb2100000000c7000415000000000000000000;                                                                          // mov
      code[ 515] = 'h0000002400000000000000eb00001500000000ea009316000000000000922100;                                                                          // moveLong
      code[ 516] = 'h00000023000000000000000000ec21000000008d000515000000000000000000;                                                                          // mov
      code[ 517] = 'h00000023000000000000000000ed2100000000c7000515000000000000000000;                                                                          // mov
      code[ 518] = 'h0000002400000000000000ed00001500000000ec009316000000000000922100;                                                                          // moveLong
      code[ 519] = 'h0000002000000000000000000000010000000000003f20000000000000000000;                                                                          // label
      code[ 520] = 'h0000002300000000000000c40002150000000000008d21000000000000000000;                                                                          // mov
      code[ 521] = 'h0000002300000000000000c70002150000000000008d21000000000000000000;                                                                          // mov
      code[ 522] = 'h00000023000000000000000000ee21000000008d000415000000000000000000;                                                                          // mov
      code[ 523] = 'h00000023000000000000000000ef2100000000ee009216000000000000000000;                                                                          // mov
      code[ 524] = 'h00000023000000000000000000f021000000008d000515000000000000000000;                                                                          // mov
      code[ 525] = 'h00000023000000000000000000f12100000000f0009216000000000000000000;                                                                          // mov
      code[ 526] = 'h00000023000000000000000000f221000000008d000415000000000000000000;                                                                          // mov
      code[ 527] = 'h0000002300000000000000f2000015000000000000ef21000000000000000000;                                                                          // mov
      code[ 528] = 'h00000023000000000000000000f321000000008d000515000000000000000000;                                                                          // mov
      code[ 529] = 'h0000002300000000000000f3000015000000000000f121000000000000000000;                                                                          // mov
      code[ 530] = 'h00000023000000000000000000f421000000008d000615000000000000000000;                                                                          // mov
      code[ 531] = 'h0000002300000000000000f4000015000000000000c421000000000000000000;                                                                          // mov
      code[ 532] = 'h00000023000000000000000000f521000000008d000615000000000000000000;                                                                          // mov
      code[ 533] = 'h0000002300000000000000f5000115000000000000c721000000000000000000;                                                                          // mov
      code[ 534] = 'h00000023000000000000008d0000150000000000000120000000000000000000;                                                                          // mov
      code[ 535] = 'h00000023000000000000000000f621000000008d000415000000000000000000;                                                                          // mov
      code[ 536] = 'h00000031000000000000000000f6210000000000000120000000000000062000;                                                                          // resize
      code[ 537] = 'h00000023000000000000000000f721000000008d000515000000000000000000;                                                                          // mov
      code[ 538] = 'h00000031000000000000000000f7210000000000000120000000000000072000;                                                                          // resize
      code[ 539] = 'h00000023000000000000000000f821000000008d000615000000000000000000;                                                                          // mov
      code[ 540] = 'h00000031000000000000000000f8210000000000000220000000000000082000;                                                                          // resize
      code[ 541] = 'h0000001f00000000000000020032210000000000000000000000000000000000;                                                                          // jmp
      code[ 542] = 'h0000001f00000000000000060034210000000000000000000000000000000000;                                                                          // jmp
      code[ 543] = 'h0000002000000000000000000000010000000000003220000000000000000000;                                                                          // label
      code[ 544] = 'h000000230000000000000000008e210000000000000120000000000000000000;                                                                          // mov
      code[ 545] = 'h0000001f00000000000000030034210000000000000000000000000000000000;                                                                          // jmp
      code[ 546] = 'h0000002000000000000000000000010000000000003320000000000000000000;                                                                          // label
      code[ 547] = 'h000000230000000000000000008e210000000000000020000000000000000000;                                                                          // mov
      code[ 548] = 'h0000002000000000000000000000010000000000003420000000000000000000;                                                                          // label
      code[ 549] = 'h0000001d00000000000000020048210000000000008e21000000000000002000;                                                                          // jNe
      code[ 550] = 'h000000230000000000000000001a210000000000008d21000000000000000000;                                                                          // mov
      code[ 551] = 'h0000002000000000000000000000010000000000004820000000000000000000;                                                                          // label
      code[ 552] = 'h0000001f00000000000000fa002d210000000000000000000000000000000000;                                                                          // jmp
      code[ 553] = 'h0000002000000000000000000000010000000000002f20000000000000000000;                                                                          // label
      code[ 554] = 'h00000023000000000000000000f921000000001a000415000000000000000000;                                                                          // mov
      code[ 555] = 'h00000005000000000000000000fa21000000000000f921000000000000042100;                                                                          // arrayIndex
      code[ 556] = 'h000000170000000000000005004921000000000000fa21000000000000002000;                                                                          // jEq
      code[ 557] = 'h0000002300000000000000060000150000000000001a21000000000000000000;                                                                          // mov
      code[ 558] = 'h0000002300000000000000060001150000000000000120000000000000000000;                                                                          // mov
      code[ 559] = 'h000000390000000000000006000215000000000000fa21000000000000012000;                                                                          // subtract
      code[ 560] = 'h0000001f00000000000000f9002a210000000000000000000000000000000000;                                                                          // jmp
      code[ 561] = 'h0000002000000000000000000000010000000000004920000000000000000000;                                                                          // label
      code[ 562] = 'h00000003000000000000000000fb21000000000000f921000000000000042100;                                                                          // arrayCountLess
      code[ 563] = 'h00000026000000000000000000fc21000000001a000615000000000000000000;                                                                          // not
      code[ 564] = 'h000000170000000000000005004a21000000000000fc21000000000000002000;                                                                          // jEq
      code[ 565] = 'h0000002300000000000000060000150000000000001a21000000000000000000;                                                                          // mov
      code[ 566] = 'h0000002300000000000000060001150000000000000020000000000000000000;                                                                          // mov
      code[ 567] = 'h000000230000000000000006000215000000000000fb21000000000000000000;                                                                          // mov
      code[ 568] = 'h0000001f00000000000000f1002a210000000000000000000000000000000000;                                                                          // jmp
      code[ 569] = 'h0000002000000000000000000000010000000000004a20000000000000000000;                                                                          // label
      code[ 570] = 'h00000023000000000000000000fd21000000001a000615000000000000000000;                                                                          // mov
      code[ 571] = 'h00000023000000000000000000fe2100000000fd00fb16000000000000000000;                                                                          // mov
      code[ 572] = 'h0000002000000000000000000000010000000000004b20000000000000000000;                                                                          // label
      code[ 573] = 'h00000023000000000000000001002100000000fe000015000000000000000000;                                                                          // mov
      code[ 574] = 'h00000023000000000000000001012100000000fe000315000000000000000000;                                                                          // mov
      code[ 575] = 'h0000002300000000000000000102210000000101000215000000000000000000;                                                                          // mov
      code[ 576] = 'h0000001c00000000000000dc004d210000000000010021000000000001022100;                                                                          // jLt
      code[ 577] = 'h0000002300000000000000000103210000000000010221000000000000000000;                                                                          // mov
      code[ 578] = 'h0000003700000000000000000103210000000000000120000000000000000000;                                                                          // shiftRight
      code[ 579] = 'h0000000000000000000000000104210000000000010321000000000000012000;                                                                          // add
      code[ 580] = 'h00000023000000000000000001052100000000fe000215000000000000000000;                                                                          // mov
      code[ 581] = 'h000000170000000000000061004f210000000000010521000000000000002000;                                                                          // jEq
      code[ 582] = 'h0000000100000000000000000106210000000000000520000000000000000000;                                                                          // array
      code[ 583] = 'h0000002300000000000001060000150000000000010321000000000000000000;                                                                          // mov
      code[ 584] = 'h0000002300000000000001060002150000000000000020000000000000000000;                                                                          // mov
      code[ 585] = 'h0000000100000000000000000107210000000000000620000000000000000000;                                                                          // array
      code[ 586] = 'h0000002300000000000001060004150000000000010721000000000000000000;                                                                          // mov
      code[ 587] = 'h0000000100000000000000000108210000000000000720000000000000000000;                                                                          // array
      code[ 588] = 'h0000002300000000000001060005150000000000010821000000000000000000;                                                                          // mov
      code[ 589] = 'h0000002300000000000001060006150000000000000020000000000000000000;                                                                          // mov
      code[ 590] = 'h0000002300000000000001060003150000000000010121000000000000000000;                                                                          // mov
      code[ 591] = 'h0000000000000000000001010001150000000101000115000000000000012000;                                                                          // add
      code[ 592] = 'h0000002300000000000001060001150000000101000115000000000000000000;                                                                          // mov
      code[ 593] = 'h00000026000000000000000001092100000000fe000615000000000000000000;                                                                          // not
      code[ 594] = 'h0000001d000000000000001d0050210000000000010921000000000000002000;                                                                          // jNe
      code[ 595] = 'h000000010000000000000000010a210000000000000820000000000000000000;                                                                          // array
      code[ 596] = 'h0000002300000000000001060006150000000000010a21000000000000000000;                                                                          // mov
      code[ 597] = 'h000000230000000000000000010b2100000000fe000415000000000000000000;                                                                          // mov
      code[ 598] = 'h000000230000000000000000010c210000000106000415000000000000000000;                                                                          // mov
      code[ 599] = 'h00000024000000000000010c000015000000010b010416000000000001032100;                                                                          // moveLong
      code[ 600] = 'h000000230000000000000000010d2100000000fe000515000000000000000000;                                                                          // mov
      code[ 601] = 'h000000230000000000000000010e210000000106000515000000000000000000;                                                                          // mov
      code[ 602] = 'h00000024000000000000010e000015000000010d010416000000000001032100;                                                                          // moveLong
      code[ 603] = 'h000000230000000000000000010f2100000000fe000615000000000000000000;                                                                          // mov
      code[ 604] = 'h0000002300000000000000000110210000000106000615000000000000000000;                                                                          // mov
      code[ 605] = 'h0000000000000000000000000111210000000000010321000000000000012000;                                                                          // add
      code[ 606] = 'h000000240000000000000110000015000000010f010416000000000001112100;                                                                          // moveLong
      code[ 607] = 'h0000002300000000000000000112210000000106000015000000000000000000;                                                                          // mov
      code[ 608] = 'h0000000000000000000000000113210000000000011221000000000000012000;                                                                          // add
      code[ 609] = 'h0000002300000000000000000114210000000106000615000000000000000000;                                                                          // mov
      code[ 610] = 'h0000002000000000000000000000010000000000005220000000000000000000;                                                                          // label
      code[ 611] = 'h0000002300000000000000000115210000000000000020000000000000000000;                                                                          // mov
      code[ 612] = 'h0000002000000000000000000000010000000000005320000000000000000000;                                                                          // label
      code[ 613] = 'h0000001900000000000000060055210000000000011521000000000001132100;                                                                          // jGe
      code[ 614] = 'h0000002300000000000000000116210000000114011516000000000000000000;                                                                          // mov
      code[ 615] = 'h0000002300000000000001160002150000000000010621000000000000000000;                                                                          // mov
      code[ 616] = 'h0000002000000000000000000000010000000000005420000000000000000000;                                                                          // label
      code[ 617] = 'h0000000000000000000000000115210000000000011521000000000000012000;                                                                          // add
      code[ 618] = 'h0000001f00000000fffffffa0053210000000000000000000000000000000000;                                                                          // jmp
      code[ 619] = 'h0000002000000000000000000000010000000000005520000000000000000000;                                                                          // label
      code[ 620] = 'h00000023000000000000000001172100000000fe000615000000000000000000;                                                                          // mov
      code[ 621] = 'h0000003100000000000000000117210000000000010421000000000000082000;                                                                          // resize
      code[ 622] = 'h0000001f00000000000000080051210000000000000000000000000000000000;                                                                          // jmp
      code[ 623] = 'h0000002000000000000000000000010000000000005020000000000000000000;                                                                          // label
      code[ 624] = 'h00000023000000000000000001182100000000fe000415000000000000000000;                                                                          // mov
      code[ 625] = 'h0000002300000000000000000119210000000106000415000000000000000000;                                                                          // mov
      code[ 626] = 'h0000002400000000000001190000150000000118010416000000000001032100;                                                                          // moveLong
      code[ 627] = 'h000000230000000000000000011a2100000000fe000515000000000000000000;                                                                          // mov
      code[ 628] = 'h000000230000000000000000011b210000000106000515000000000000000000;                                                                          // mov
      code[ 629] = 'h00000024000000000000011b000015000000011a010416000000000001032100;                                                                          // moveLong
      code[ 630] = 'h0000002000000000000000000000010000000000005120000000000000000000;                                                                          // label
      code[ 631] = 'h0000002300000000000000fe0000150000000000010321000000000000000000;                                                                          // mov
      code[ 632] = 'h0000002300000000000001060002150000000000010521000000000000000000;                                                                          // mov
      code[ 633] = 'h000000230000000000000000011c210000000105000015000000000000000000;                                                                          // mov
      code[ 634] = 'h000000230000000000000000011d210000000105000615000000000000000000;                                                                          // mov
      code[ 635] = 'h000000230000000000000000011e21000000011d011c16000000000000000000;                                                                          // mov
      code[ 636] = 'h0000001d00000000000000130056210000000000011e21000000000000fe2100;                                                                          // jNe
      code[ 637] = 'h000000230000000000000000011f2100000000fe000415000000000000000000;                                                                          // mov
      code[ 638] = 'h000000230000000000000000012021000000011f010316000000000000000000;                                                                          // mov
      code[ 639] = 'h0000002300000000000000000121210000000105000415000000000000000000;                                                                          // mov
      code[ 640] = 'h000000230000000000000121011c160000000000012021000000000000000000;                                                                          // mov
      code[ 641] = 'h00000023000000000000000001222100000000fe000515000000000000000000;                                                                          // mov
      code[ 642] = 'h0000002300000000000000000123210000000122010316000000000000000000;                                                                          // mov
      code[ 643] = 'h0000002300000000000000000124210000000105000515000000000000000000;                                                                          // mov
      code[ 644] = 'h000000230000000000000124011c160000000000012321000000000000000000;                                                                          // mov
      code[ 645] = 'h00000023000000000000000001252100000000fe000415000000000000000000;                                                                          // mov
      code[ 646] = 'h0000003100000000000000000125210000000000010321000000000000062000;                                                                          // resize
      code[ 647] = 'h00000023000000000000000001262100000000fe000515000000000000000000;                                                                          // mov
      code[ 648] = 'h0000003100000000000000000126210000000000010321000000000000072000;                                                                          // resize
      code[ 649] = 'h0000000000000000000000000127210000000000011c21000000000000012000;                                                                          // add
      code[ 650] = 'h0000002300000000000001050000150000000000012721000000000000000000;                                                                          // mov
      code[ 651] = 'h0000002300000000000000000128210000000105000615000000000000000000;                                                                          // mov
      code[ 652] = 'h0000002300000000000001280127160000000000010621000000000000000000;                                                                          // mov
      code[ 653] = 'h0000001f000000000000008c004c210000000000000000000000000000000000;                                                                          // jmp
      code[ 654] = 'h0000001f00000000000000170057210000000000000000000000000000000000;                                                                          // jmp
      code[ 655] = 'h0000002000000000000000000000010000000000005620000000000000000000;                                                                          // label
      code[ 656] = 'h0000000f00000000000000000000010000000000010521000000000000002000;                                                                          // assertNe
      code[ 657] = 'h0000002300000000000000000129210000000105000615000000000000000000;                                                                          // mov
      code[ 658] = 'h000000050000000000000000012a210000000000012921000000000000fe2100;                                                                          // arrayIndex
      code[ 659] = 'h000000390000000000000000012a210000000000012a21000000000000012000;                                                                          // subtract
      code[ 660] = 'h000000230000000000000000012b2100000000fe000415000000000000000000;                                                                          // mov
      code[ 661] = 'h000000230000000000000000012c21000000012b010316000000000000000000;                                                                          // mov
      code[ 662] = 'h000000230000000000000000012d2100000000fe000515000000000000000000;                                                                          // mov
      code[ 663] = 'h000000230000000000000000012e21000000012d010316000000000000000000;                                                                          // mov
      code[ 664] = 'h000000230000000000000000012f2100000000fe000415000000000000000000;                                                                          // mov
      code[ 665] = 'h000000310000000000000000012f210000000000010321000000000000062000;                                                                          // resize
      code[ 666] = 'h00000023000000000000000001302100000000fe000515000000000000000000;                                                                          // mov
      code[ 667] = 'h0000003100000000000000000130210000000000010321000000000000072000;                                                                          // resize
      code[ 668] = 'h0000002300000000000000000131210000000105000415000000000000000000;                                                                          // mov
      code[ 669] = 'h000000380000000000000131012a160000000000012c21000000000000000000;                                                                          // shiftUp
      code[ 670] = 'h0000002300000000000000000132210000000105000515000000000000000000;                                                                          // mov
      code[ 671] = 'h000000380000000000000132012a160000000000012e21000000000000000000;                                                                          // shiftUp
      code[ 672] = 'h0000002300000000000000000133210000000105000615000000000000000000;                                                                          // mov
      code[ 673] = 'h0000000000000000000000000134210000000000012a21000000000000012000;                                                                          // add
      code[ 674] = 'h0000003800000000000001330134160000000000010621000000000000000000;                                                                          // shiftUp
      code[ 675] = 'h0000000000000000000001050000150000000105000015000000000000012000;                                                                          // add
      code[ 676] = 'h0000001f0000000000000075004c210000000000000000000000000000000000;                                                                          // jmp
      code[ 677] = 'h0000002000000000000000000000010000000000005720000000000000000000;                                                                          // label
      code[ 678] = 'h0000002000000000000000000000010000000000004f20000000000000000000;                                                                          // label
      code[ 679] = 'h0000000100000000000000000135210000000000000520000000000000000000;                                                                          // array
      code[ 680] = 'h0000002300000000000001350000150000000000010321000000000000000000;                                                                          // mov
      code[ 681] = 'h0000002300000000000001350002150000000000000020000000000000000000;                                                                          // mov
      code[ 682] = 'h0000000100000000000000000136210000000000000620000000000000000000;                                                                          // array
      code[ 683] = 'h0000002300000000000001350004150000000000013621000000000000000000;                                                                          // mov
      code[ 684] = 'h0000000100000000000000000137210000000000000720000000000000000000;                                                                          // array
      code[ 685] = 'h0000002300000000000001350005150000000000013721000000000000000000;                                                                          // mov
      code[ 686] = 'h0000002300000000000001350006150000000000000020000000000000000000;                                                                          // mov
      code[ 687] = 'h0000002300000000000001350003150000000000010121000000000000000000;                                                                          // mov
      code[ 688] = 'h0000000000000000000001010001150000000101000115000000000000012000;                                                                          // add
      code[ 689] = 'h0000002300000000000001350001150000000101000115000000000000000000;                                                                          // mov
      code[ 690] = 'h0000000100000000000000000138210000000000000520000000000000000000;                                                                          // array
      code[ 691] = 'h0000002300000000000001380000150000000000010321000000000000000000;                                                                          // mov
      code[ 692] = 'h0000002300000000000001380002150000000000000020000000000000000000;                                                                          // mov
      code[ 693] = 'h0000000100000000000000000139210000000000000620000000000000000000;                                                                          // array
      code[ 694] = 'h0000002300000000000001380004150000000000013921000000000000000000;                                                                          // mov
      code[ 695] = 'h000000010000000000000000013a210000000000000720000000000000000000;                                                                          // array
      code[ 696] = 'h0000002300000000000001380005150000000000013a21000000000000000000;                                                                          // mov
      code[ 697] = 'h0000002300000000000001380006150000000000000020000000000000000000;                                                                          // mov
      code[ 698] = 'h0000002300000000000001380003150000000000010121000000000000000000;                                                                          // mov
      code[ 699] = 'h0000000000000000000001010001150000000101000115000000000000012000;                                                                          // add
      code[ 700] = 'h0000002300000000000001380001150000000101000115000000000000000000;                                                                          // mov
      code[ 701] = 'h000000260000000000000000013b2100000000fe000615000000000000000000;                                                                          // not
      code[ 702] = 'h0000001d00000000000000340058210000000000013b21000000000000002000;                                                                          // jNe
      code[ 703] = 'h000000010000000000000000013c210000000000000820000000000000000000;                                                                          // array
      code[ 704] = 'h0000002300000000000001350006150000000000013c21000000000000000000;                                                                          // mov
      code[ 705] = 'h000000010000000000000000013d210000000000000820000000000000000000;                                                                          // array
      code[ 706] = 'h0000002300000000000001380006150000000000013d21000000000000000000;                                                                          // mov
      code[ 707] = 'h000000230000000000000000013e2100000000fe000415000000000000000000;                                                                          // mov
      code[ 708] = 'h000000230000000000000000013f210000000135000415000000000000000000;                                                                          // mov
      code[ 709] = 'h00000024000000000000013f000015000000013e000015000000000001032100;                                                                          // moveLong
      code[ 710] = 'h00000023000000000000000001402100000000fe000515000000000000000000;                                                                          // mov
      code[ 711] = 'h0000002300000000000000000141210000000135000515000000000000000000;                                                                          // mov
      code[ 712] = 'h0000002400000000000001410000150000000140000015000000000001032100;                                                                          // moveLong
      code[ 713] = 'h00000023000000000000000001422100000000fe000615000000000000000000;                                                                          // mov
      code[ 714] = 'h0000002300000000000000000143210000000135000615000000000000000000;                                                                          // mov
      code[ 715] = 'h0000000000000000000000000144210000000000010321000000000000012000;                                                                          // add
      code[ 716] = 'h0000002400000000000001430000150000000142000015000000000001442100;                                                                          // moveLong
      code[ 717] = 'h00000023000000000000000001452100000000fe000415000000000000000000;                                                                          // mov
      code[ 718] = 'h0000002300000000000000000146210000000138000415000000000000000000;                                                                          // mov
      code[ 719] = 'h0000002400000000000001460000150000000145010416000000000001032100;                                                                          // moveLong
      code[ 720] = 'h00000023000000000000000001472100000000fe000515000000000000000000;                                                                          // mov
      code[ 721] = 'h0000002300000000000000000148210000000138000515000000000000000000;                                                                          // mov
      code[ 722] = 'h0000002400000000000001480000150000000147010416000000000001032100;                                                                          // moveLong
      code[ 723] = 'h00000023000000000000000001492100000000fe000615000000000000000000;                                                                          // mov
      code[ 724] = 'h000000230000000000000000014a210000000138000615000000000000000000;                                                                          // mov
      code[ 725] = 'h000000000000000000000000014b210000000000010321000000000000012000;                                                                          // add
      code[ 726] = 'h00000024000000000000014a00001500000001490104160000000000014b2100;                                                                          // moveLong
      code[ 727] = 'h000000230000000000000000014c210000000135000015000000000000000000;                                                                          // mov
      code[ 728] = 'h000000000000000000000000014d210000000000014c21000000000000012000;                                                                          // add
      code[ 729] = 'h000000230000000000000000014e210000000135000615000000000000000000;                                                                          // mov
      code[ 730] = 'h0000002000000000000000000000010000000000005a20000000000000000000;                                                                          // label
      code[ 731] = 'h000000230000000000000000014f210000000000000020000000000000000000;                                                                          // mov
      code[ 732] = 'h0000002000000000000000000000010000000000005b20000000000000000000;                                                                          // label
      code[ 733] = 'h000000190000000000000006005d210000000000014f210000000000014d2100;                                                                          // jGe
      code[ 734] = 'h000000230000000000000000015021000000014e014f16000000000000000000;                                                                          // mov
      code[ 735] = 'h0000002300000000000001500002150000000000013521000000000000000000;                                                                          // mov
      code[ 736] = 'h0000002000000000000000000000010000000000005c20000000000000000000;                                                                          // label
      code[ 737] = 'h000000000000000000000000014f210000000000014f21000000000000012000;                                                                          // add
      code[ 738] = 'h0000001f00000000fffffffa005b210000000000000000000000000000000000;                                                                          // jmp
      code[ 739] = 'h0000002000000000000000000000010000000000005d20000000000000000000;                                                                          // label
      code[ 740] = 'h0000002300000000000000000151210000000138000015000000000000000000;                                                                          // mov
      code[ 741] = 'h0000000000000000000000000152210000000000015121000000000000012000;                                                                          // add
      code[ 742] = 'h0000002300000000000000000153210000000138000615000000000000000000;                                                                          // mov
      code[ 743] = 'h0000002000000000000000000000010000000000005e20000000000000000000;                                                                          // label
      code[ 744] = 'h0000002300000000000000000154210000000000000020000000000000000000;                                                                          // mov
      code[ 745] = 'h0000002000000000000000000000010000000000005f20000000000000000000;                                                                          // label
      code[ 746] = 'h0000001900000000000000060061210000000000015421000000000001522100;                                                                          // jGe
      code[ 747] = 'h0000002300000000000000000155210000000153015416000000000000000000;                                                                          // mov
      code[ 748] = 'h0000002300000000000001550002150000000000013821000000000000000000;                                                                          // mov
      code[ 749] = 'h0000002000000000000000000000010000000000006020000000000000000000;                                                                          // label
      code[ 750] = 'h0000000000000000000000000154210000000000015421000000000000012000;                                                                          // add
      code[ 751] = 'h0000001f00000000fffffffa005f210000000000000000000000000000000000;                                                                          // jmp
      code[ 752] = 'h0000002000000000000000000000010000000000006120000000000000000000;                                                                          // label
      code[ 753] = 'h0000001f00000000000000100059210000000000000000000000000000000000;                                                                          // jmp
      code[ 754] = 'h0000002000000000000000000000010000000000005820000000000000000000;                                                                          // label
      code[ 755] = 'h0000000100000000000000000156210000000000000820000000000000000000;                                                                          // array
      code[ 756] = 'h0000002300000000000000fe0006150000000000015621000000000000000000;                                                                          // mov
      code[ 757] = 'h00000023000000000000000001572100000000fe000415000000000000000000;                                                                          // mov
      code[ 758] = 'h0000002300000000000000000158210000000135000415000000000000000000;                                                                          // mov
      code[ 759] = 'h0000002400000000000001580000150000000157000015000000000001032100;                                                                          // moveLong
      code[ 760] = 'h00000023000000000000000001592100000000fe000515000000000000000000;                                                                          // mov
      code[ 761] = 'h000000230000000000000000015a210000000135000515000000000000000000;                                                                          // mov
      code[ 762] = 'h00000024000000000000015a0000150000000159000015000000000001032100;                                                                          // moveLong
      code[ 763] = 'h000000230000000000000000015b2100000000fe000415000000000000000000;                                                                          // mov
      code[ 764] = 'h000000230000000000000000015c210000000138000415000000000000000000;                                                                          // mov
      code[ 765] = 'h00000024000000000000015c000015000000015b010416000000000001032100;                                                                          // moveLong
      code[ 766] = 'h000000230000000000000000015d2100000000fe000515000000000000000000;                                                                          // mov
      code[ 767] = 'h000000230000000000000000015e210000000138000515000000000000000000;                                                                          // mov
      code[ 768] = 'h00000024000000000000015e000015000000015d010416000000000001032100;                                                                          // moveLong
      code[ 769] = 'h0000002000000000000000000000010000000000005920000000000000000000;                                                                          // label
      code[ 770] = 'h000000230000000000000135000215000000000000fe21000000000000000000;                                                                          // mov
      code[ 771] = 'h000000230000000000000138000215000000000000fe21000000000000000000;                                                                          // mov
      code[ 772] = 'h000000230000000000000000015f2100000000fe000415000000000000000000;                                                                          // mov
      code[ 773] = 'h000000230000000000000000016021000000015f010316000000000000000000;                                                                          // mov
      code[ 774] = 'h00000023000000000000000001612100000000fe000515000000000000000000;                                                                          // mov
      code[ 775] = 'h0000002300000000000000000162210000000161010316000000000000000000;                                                                          // mov
      code[ 776] = 'h00000023000000000000000001632100000000fe000415000000000000000000;                                                                          // mov
      code[ 777] = 'h0000002300000000000001630000150000000000016021000000000000000000;                                                                          // mov
      code[ 778] = 'h00000023000000000000000001642100000000fe000515000000000000000000;                                                                          // mov
      code[ 779] = 'h0000002300000000000001640000150000000000016221000000000000000000;                                                                          // mov
      code[ 780] = 'h00000023000000000000000001652100000000fe000615000000000000000000;                                                                          // mov
      code[ 781] = 'h0000002300000000000001650000150000000000013521000000000000000000;                                                                          // mov
      code[ 782] = 'h00000023000000000000000001662100000000fe000615000000000000000000;                                                                          // mov
      code[ 783] = 'h0000002300000000000001660001150000000000013821000000000000000000;                                                                          // mov
      code[ 784] = 'h0000002300000000000000fe0000150000000000000120000000000000000000;                                                                          // mov
      code[ 785] = 'h00000023000000000000000001672100000000fe000415000000000000000000;                                                                          // mov
      code[ 786] = 'h0000003100000000000000000167210000000000000120000000000000062000;                                                                          // resize
      code[ 787] = 'h00000023000000000000000001682100000000fe000515000000000000000000;                                                                          // mov
      code[ 788] = 'h0000003100000000000000000168210000000000000120000000000000072000;                                                                          // resize
      code[ 789] = 'h00000023000000000000000001692100000000fe000615000000000000000000;                                                                          // mov
      code[ 790] = 'h0000003100000000000000000169210000000000000220000000000000082000;                                                                          // resize
      code[ 791] = 'h0000001f0000000000000002004c210000000000000000000000000000000000;                                                                          // jmp
      code[ 792] = 'h0000001f0000000000000006004e210000000000000000000000000000000000;                                                                          // jmp
      code[ 793] = 'h0000002000000000000000000000010000000000004c20000000000000000000;                                                                          // label
      code[ 794] = 'h00000023000000000000000000ff210000000000000120000000000000000000;                                                                          // mov
      code[ 795] = 'h0000001f0000000000000003004e210000000000000000000000000000000000;                                                                          // jmp
      code[ 796] = 'h0000002000000000000000000000010000000000004d20000000000000000000;                                                                          // label
      code[ 797] = 'h00000023000000000000000000ff210000000000000020000000000000000000;                                                                          // mov
      code[ 798] = 'h0000002000000000000000000000010000000000004e20000000000000000000;                                                                          // label
      code[ 799] = 'h0000001d0000000000000002006221000000000000ff21000000000000002000;                                                                          // jNe
      code[ 800] = 'h000000230000000000000000001a21000000000000fe21000000000000000000;                                                                          // mov
      code[ 801] = 'h0000002000000000000000000000010000000000006220000000000000000000;                                                                          // label
      code[ 802] = 'h0000002000000000000000000000010000000000002d20000000000000000000;                                                                          // label
      code[ 803] = 'h0000000000000000000000000086210000000000008621000000000000012000;                                                                          // add
      code[ 804] = 'h0000001f00000000fffffe0e002c210000000000000000000000000000000000;                                                                          // jmp
      code[ 805] = 'h0000002000000000000000000000010000000000002e20000000000000000000;                                                                          // label
      code[ 806] = 'h0000000800000000000000000000010000000000000000000000000000000000;                                                                          // assert
      code[ 807] = 'h0000002000000000000000000000010000000000002820000000000000000000;                                                                          // label
      code[ 808] = 'h0000002000000000000000000000010000000000002920000000000000000000;                                                                          // label
      code[ 809] = 'h0000002000000000000000000000010000000000002a20000000000000000000;                                                                          // label
      code[ 810] = 'h000000230000000000000000016a210000000006000015000000000000000000;                                                                          // mov
      code[ 811] = 'h000000230000000000000000016b210000000006000115000000000000000000;                                                                          // mov
      code[ 812] = 'h000000230000000000000000016c210000000006000215000000000000000000;                                                                          // mov
      code[ 813] = 'h0000001d00000000000000040063210000000000016b21000000000000012000;                                                                          // jNe
      code[ 814] = 'h000000230000000000000000016d21000000016a000515000000000000000000;                                                                          // mov
      code[ 815] = 'h00000023000000000000016d016c160000000000000521000000000000000000;                                                                          // mov
      code[ 816] = 'h0000001f00000000000000f70009210000000000000000000000000000000000;                                                                          // jmp
      code[ 817] = 'h0000002000000000000000000000010000000000006320000000000000000000;                                                                          // label
      code[ 818] = 'h0000001d00000000000000080064210000000000016b21000000000000022000;                                                                          // jNe
      code[ 819] = 'h000000000000000000000000016e210000000000016c21000000000000012000;                                                                          // add
      code[ 820] = 'h000000230000000000000000016f21000000016a000415000000000000000000;                                                                          // mov
      code[ 821] = 'h00000038000000000000016f016e160000000000000421000000000000000000;                                                                          // shiftUp
      code[ 822] = 'h000000230000000000000000017021000000016a000515000000000000000000;                                                                          // mov
      code[ 823] = 'h000000380000000000000170016e160000000000000521000000000000000000;                                                                          // shiftUp
      code[ 824] = 'h00000000000000000000016a000015000000016a000015000000000000012000;                                                                          // add
      code[ 825] = 'h0000001f00000000000000070065210000000000000000000000000000000000;                                                                          // jmp
      code[ 826] = 'h0000002000000000000000000000010000000000006420000000000000000000;                                                                          // label
      code[ 827] = 'h000000230000000000000000017121000000016a000415000000000000000000;                                                                          // mov
      code[ 828] = 'h000000380000000000000171016c160000000000000421000000000000000000;                                                                          // shiftUp
      code[ 829] = 'h000000230000000000000000017221000000016a000515000000000000000000;                                                                          // mov
      code[ 830] = 'h000000380000000000000172016c160000000000000521000000000000000000;                                                                          // shiftUp
      code[ 831] = 'h00000000000000000000016a000015000000016a000015000000000000012000;                                                                          // add
      code[ 832] = 'h0000002000000000000000000000010000000000006520000000000000000000;                                                                          // label
      code[ 833] = 'h0000000000000000000000030000150000000003000015000000000000012000;                                                                          // add
      code[ 834] = 'h0000002000000000000000000000010000000000006620000000000000000000;                                                                          // label
      code[ 835] = 'h000000230000000000000000017421000000016a000015000000000000000000;                                                                          // mov
      code[ 836] = 'h000000230000000000000000017521000000016a000315000000000000000000;                                                                          // mov
      code[ 837] = 'h0000002300000000000000000176210000000175000215000000000000000000;                                                                          // mov
      code[ 838] = 'h0000001c00000000000000dc0068210000000000017421000000000001762100;                                                                          // jLt
      code[ 839] = 'h0000002300000000000000000177210000000000017621000000000000000000;                                                                          // mov
      code[ 840] = 'h0000003700000000000000000177210000000000000120000000000000000000;                                                                          // shiftRight
      code[ 841] = 'h0000000000000000000000000178210000000000017721000000000000012000;                                                                          // add
      code[ 842] = 'h000000230000000000000000017921000000016a000215000000000000000000;                                                                          // mov
      code[ 843] = 'h000000170000000000000061006a210000000000017921000000000000002000;                                                                          // jEq
      code[ 844] = 'h000000010000000000000000017a210000000000000520000000000000000000;                                                                          // array
      code[ 845] = 'h00000023000000000000017a0000150000000000017721000000000000000000;                                                                          // mov
      code[ 846] = 'h00000023000000000000017a0002150000000000000020000000000000000000;                                                                          // mov
      code[ 847] = 'h000000010000000000000000017b210000000000000620000000000000000000;                                                                          // array
      code[ 848] = 'h00000023000000000000017a0004150000000000017b21000000000000000000;                                                                          // mov
      code[ 849] = 'h000000010000000000000000017c210000000000000720000000000000000000;                                                                          // array
      code[ 850] = 'h00000023000000000000017a0005150000000000017c21000000000000000000;                                                                          // mov
      code[ 851] = 'h00000023000000000000017a0006150000000000000020000000000000000000;                                                                          // mov
      code[ 852] = 'h00000023000000000000017a0003150000000000017521000000000000000000;                                                                          // mov
      code[ 853] = 'h0000000000000000000001750001150000000175000115000000000000012000;                                                                          // add
      code[ 854] = 'h00000023000000000000017a0001150000000175000115000000000000000000;                                                                          // mov
      code[ 855] = 'h000000260000000000000000017d21000000016a000615000000000000000000;                                                                          // not
      code[ 856] = 'h0000001d000000000000001d006b210000000000017d21000000000000002000;                                                                          // jNe
      code[ 857] = 'h000000010000000000000000017e210000000000000820000000000000000000;                                                                          // array
      code[ 858] = 'h00000023000000000000017a0006150000000000017e21000000000000000000;                                                                          // mov
      code[ 859] = 'h000000230000000000000000017f21000000016a000415000000000000000000;                                                                          // mov
      code[ 860] = 'h000000230000000000000000018021000000017a000415000000000000000000;                                                                          // mov
      code[ 861] = 'h000000240000000000000180000015000000017f017816000000000001772100;                                                                          // moveLong
      code[ 862] = 'h000000230000000000000000018121000000016a000515000000000000000000;                                                                          // mov
      code[ 863] = 'h000000230000000000000000018221000000017a000515000000000000000000;                                                                          // mov
      code[ 864] = 'h0000002400000000000001820000150000000181017816000000000001772100;                                                                          // moveLong
      code[ 865] = 'h000000230000000000000000018321000000016a000615000000000000000000;                                                                          // mov
      code[ 866] = 'h000000230000000000000000018421000000017a000615000000000000000000;                                                                          // mov
      code[ 867] = 'h0000000000000000000000000185210000000000017721000000000000012000;                                                                          // add
      code[ 868] = 'h0000002400000000000001840000150000000183017816000000000001852100;                                                                          // moveLong
      code[ 869] = 'h000000230000000000000000018621000000017a000015000000000000000000;                                                                          // mov
      code[ 870] = 'h0000000000000000000000000187210000000000018621000000000000012000;                                                                          // add
      code[ 871] = 'h000000230000000000000000018821000000017a000615000000000000000000;                                                                          // mov
      code[ 872] = 'h0000002000000000000000000000010000000000006d20000000000000000000;                                                                          // label
      code[ 873] = 'h0000002300000000000000000189210000000000000020000000000000000000;                                                                          // mov
      code[ 874] = 'h0000002000000000000000000000010000000000006e20000000000000000000;                                                                          // label
      code[ 875] = 'h0000001900000000000000060070210000000000018921000000000001872100;                                                                          // jGe
      code[ 876] = 'h000000230000000000000000018a210000000188018916000000000000000000;                                                                          // mov
      code[ 877] = 'h00000023000000000000018a0002150000000000017a21000000000000000000;                                                                          // mov
      code[ 878] = 'h0000002000000000000000000000010000000000006f20000000000000000000;                                                                          // label
      code[ 879] = 'h0000000000000000000000000189210000000000018921000000000000012000;                                                                          // add
      code[ 880] = 'h0000001f00000000fffffffa006e210000000000000000000000000000000000;                                                                          // jmp
      code[ 881] = 'h0000002000000000000000000000010000000000007020000000000000000000;                                                                          // label
      code[ 882] = 'h000000230000000000000000018b21000000016a000615000000000000000000;                                                                          // mov
      code[ 883] = 'h000000310000000000000000018b210000000000017821000000000000082000;                                                                          // resize
      code[ 884] = 'h0000001f0000000000000008006c210000000000000000000000000000000000;                                                                          // jmp
      code[ 885] = 'h0000002000000000000000000000010000000000006b20000000000000000000;                                                                          // label
      code[ 886] = 'h000000230000000000000000018c21000000016a000415000000000000000000;                                                                          // mov
      code[ 887] = 'h000000230000000000000000018d21000000017a000415000000000000000000;                                                                          // mov
      code[ 888] = 'h00000024000000000000018d000015000000018c017816000000000001772100;                                                                          // moveLong
      code[ 889] = 'h000000230000000000000000018e21000000016a000515000000000000000000;                                                                          // mov
      code[ 890] = 'h000000230000000000000000018f21000000017a000515000000000000000000;                                                                          // mov
      code[ 891] = 'h00000024000000000000018f000015000000018e017816000000000001772100;                                                                          // moveLong
      code[ 892] = 'h0000002000000000000000000000010000000000006c20000000000000000000;                                                                          // label
      code[ 893] = 'h00000023000000000000016a0000150000000000017721000000000000000000;                                                                          // mov
      code[ 894] = 'h00000023000000000000017a0002150000000000017921000000000000000000;                                                                          // mov
      code[ 895] = 'h0000002300000000000000000190210000000179000015000000000000000000;                                                                          // mov
      code[ 896] = 'h0000002300000000000000000191210000000179000615000000000000000000;                                                                          // mov
      code[ 897] = 'h0000002300000000000000000192210000000191019016000000000000000000;                                                                          // mov
      code[ 898] = 'h0000001d000000000000001300712100000000000192210000000000016a2100;                                                                          // jNe
      code[ 899] = 'h000000230000000000000000019321000000016a000415000000000000000000;                                                                          // mov
      code[ 900] = 'h0000002300000000000000000194210000000193017716000000000000000000;                                                                          // mov
      code[ 901] = 'h0000002300000000000000000195210000000179000415000000000000000000;                                                                          // mov
      code[ 902] = 'h0000002300000000000001950190160000000000019421000000000000000000;                                                                          // mov
      code[ 903] = 'h000000230000000000000000019621000000016a000515000000000000000000;                                                                          // mov
      code[ 904] = 'h0000002300000000000000000197210000000196017716000000000000000000;                                                                          // mov
      code[ 905] = 'h0000002300000000000000000198210000000179000515000000000000000000;                                                                          // mov
      code[ 906] = 'h0000002300000000000001980190160000000000019721000000000000000000;                                                                          // mov
      code[ 907] = 'h000000230000000000000000019921000000016a000415000000000000000000;                                                                          // mov
      code[ 908] = 'h0000003100000000000000000199210000000000017721000000000000062000;                                                                          // resize
      code[ 909] = 'h000000230000000000000000019a21000000016a000515000000000000000000;                                                                          // mov
      code[ 910] = 'h000000310000000000000000019a210000000000017721000000000000072000;                                                                          // resize
      code[ 911] = 'h000000000000000000000000019b210000000000019021000000000000012000;                                                                          // add
      code[ 912] = 'h0000002300000000000001790000150000000000019b21000000000000000000;                                                                          // mov
      code[ 913] = 'h000000230000000000000000019c210000000179000615000000000000000000;                                                                          // mov
      code[ 914] = 'h00000023000000000000019c019b160000000000017a21000000000000000000;                                                                          // mov
      code[ 915] = 'h0000001f000000000000008c0067210000000000000000000000000000000000;                                                                          // jmp
      code[ 916] = 'h0000001f00000000000000170072210000000000000000000000000000000000;                                                                          // jmp
      code[ 917] = 'h0000002000000000000000000000010000000000007120000000000000000000;                                                                          // label
      code[ 918] = 'h0000000f00000000000000000000010000000000017921000000000000002000;                                                                          // assertNe
      code[ 919] = 'h000000230000000000000000019d210000000179000615000000000000000000;                                                                          // mov
      code[ 920] = 'h000000050000000000000000019e210000000000019d210000000000016a2100;                                                                          // arrayIndex
      code[ 921] = 'h000000390000000000000000019e210000000000019e21000000000000012000;                                                                          // subtract
      code[ 922] = 'h000000230000000000000000019f21000000016a000415000000000000000000;                                                                          // mov
      code[ 923] = 'h00000023000000000000000001a021000000019f017716000000000000000000;                                                                          // mov
      code[ 924] = 'h00000023000000000000000001a121000000016a000515000000000000000000;                                                                          // mov
      code[ 925] = 'h00000023000000000000000001a22100000001a1017716000000000000000000;                                                                          // mov
      code[ 926] = 'h00000023000000000000000001a321000000016a000415000000000000000000;                                                                          // mov
      code[ 927] = 'h00000031000000000000000001a3210000000000017721000000000000062000;                                                                          // resize
      code[ 928] = 'h00000023000000000000000001a421000000016a000515000000000000000000;                                                                          // mov
      code[ 929] = 'h00000031000000000000000001a4210000000000017721000000000000072000;                                                                          // resize
      code[ 930] = 'h00000023000000000000000001a5210000000179000415000000000000000000;                                                                          // mov
      code[ 931] = 'h0000003800000000000001a5019e16000000000001a021000000000000000000;                                                                          // shiftUp
      code[ 932] = 'h00000023000000000000000001a6210000000179000515000000000000000000;                                                                          // mov
      code[ 933] = 'h0000003800000000000001a6019e16000000000001a221000000000000000000;                                                                          // shiftUp
      code[ 934] = 'h00000023000000000000000001a7210000000179000615000000000000000000;                                                                          // mov
      code[ 935] = 'h00000000000000000000000001a8210000000000019e21000000000000012000;                                                                          // add
      code[ 936] = 'h0000003800000000000001a701a8160000000000017a21000000000000000000;                                                                          // shiftUp
      code[ 937] = 'h0000000000000000000001790000150000000179000015000000000000012000;                                                                          // add
      code[ 938] = 'h0000001f00000000000000750067210000000000000000000000000000000000;                                                                          // jmp
      code[ 939] = 'h0000002000000000000000000000010000000000007220000000000000000000;                                                                          // label
      code[ 940] = 'h0000002000000000000000000000010000000000006a20000000000000000000;                                                                          // label
      code[ 941] = 'h00000001000000000000000001a9210000000000000520000000000000000000;                                                                          // array
      code[ 942] = 'h0000002300000000000001a90000150000000000017721000000000000000000;                                                                          // mov
      code[ 943] = 'h0000002300000000000001a90002150000000000000020000000000000000000;                                                                          // mov
      code[ 944] = 'h00000001000000000000000001aa210000000000000620000000000000000000;                                                                          // array
      code[ 945] = 'h0000002300000000000001a9000415000000000001aa21000000000000000000;                                                                          // mov
      code[ 946] = 'h00000001000000000000000001ab210000000000000720000000000000000000;                                                                          // array
      code[ 947] = 'h0000002300000000000001a9000515000000000001ab21000000000000000000;                                                                          // mov
      code[ 948] = 'h0000002300000000000001a90006150000000000000020000000000000000000;                                                                          // mov
      code[ 949] = 'h0000002300000000000001a90003150000000000017521000000000000000000;                                                                          // mov
      code[ 950] = 'h0000000000000000000001750001150000000175000115000000000000012000;                                                                          // add
      code[ 951] = 'h0000002300000000000001a90001150000000175000115000000000000000000;                                                                          // mov
      code[ 952] = 'h00000001000000000000000001ac210000000000000520000000000000000000;                                                                          // array
      code[ 953] = 'h0000002300000000000001ac0000150000000000017721000000000000000000;                                                                          // mov
      code[ 954] = 'h0000002300000000000001ac0002150000000000000020000000000000000000;                                                                          // mov
      code[ 955] = 'h00000001000000000000000001ad210000000000000620000000000000000000;                                                                          // array
      code[ 956] = 'h0000002300000000000001ac000415000000000001ad21000000000000000000;                                                                          // mov
      code[ 957] = 'h00000001000000000000000001ae210000000000000720000000000000000000;                                                                          // array
      code[ 958] = 'h0000002300000000000001ac000515000000000001ae21000000000000000000;                                                                          // mov
      code[ 959] = 'h0000002300000000000001ac0006150000000000000020000000000000000000;                                                                          // mov
      code[ 960] = 'h0000002300000000000001ac0003150000000000017521000000000000000000;                                                                          // mov
      code[ 961] = 'h0000000000000000000001750001150000000175000115000000000000012000;                                                                          // add
      code[ 962] = 'h0000002300000000000001ac0001150000000175000115000000000000000000;                                                                          // mov
      code[ 963] = 'h00000026000000000000000001af21000000016a000615000000000000000000;                                                                          // not
      code[ 964] = 'h0000001d0000000000000034007321000000000001af21000000000000002000;                                                                          // jNe
      code[ 965] = 'h00000001000000000000000001b0210000000000000820000000000000000000;                                                                          // array
      code[ 966] = 'h0000002300000000000001a9000615000000000001b021000000000000000000;                                                                          // mov
      code[ 967] = 'h00000001000000000000000001b1210000000000000820000000000000000000;                                                                          // array
      code[ 968] = 'h0000002300000000000001ac000615000000000001b121000000000000000000;                                                                          // mov
      code[ 969] = 'h00000023000000000000000001b221000000016a000415000000000000000000;                                                                          // mov
      code[ 970] = 'h00000023000000000000000001b32100000001a9000415000000000000000000;                                                                          // mov
      code[ 971] = 'h0000002400000000000001b300001500000001b2000015000000000001772100;                                                                          // moveLong
      code[ 972] = 'h00000023000000000000000001b421000000016a000515000000000000000000;                                                                          // mov
      code[ 973] = 'h00000023000000000000000001b52100000001a9000515000000000000000000;                                                                          // mov
      code[ 974] = 'h0000002400000000000001b500001500000001b4000015000000000001772100;                                                                          // moveLong
      code[ 975] = 'h00000023000000000000000001b621000000016a000615000000000000000000;                                                                          // mov
      code[ 976] = 'h00000023000000000000000001b72100000001a9000615000000000000000000;                                                                          // mov
      code[ 977] = 'h00000000000000000000000001b8210000000000017721000000000000012000;                                                                          // add
      code[ 978] = 'h0000002400000000000001b700001500000001b6000015000000000001b82100;                                                                          // moveLong
      code[ 979] = 'h00000023000000000000000001b921000000016a000415000000000000000000;                                                                          // mov
      code[ 980] = 'h00000023000000000000000001ba2100000001ac000415000000000000000000;                                                                          // mov
      code[ 981] = 'h0000002400000000000001ba00001500000001b9017816000000000001772100;                                                                          // moveLong
      code[ 982] = 'h00000023000000000000000001bb21000000016a000515000000000000000000;                                                                          // mov
      code[ 983] = 'h00000023000000000000000001bc2100000001ac000515000000000000000000;                                                                          // mov
      code[ 984] = 'h0000002400000000000001bc00001500000001bb017816000000000001772100;                                                                          // moveLong
      code[ 985] = 'h00000023000000000000000001bd21000000016a000615000000000000000000;                                                                          // mov
      code[ 986] = 'h00000023000000000000000001be2100000001ac000615000000000000000000;                                                                          // mov
      code[ 987] = 'h00000000000000000000000001bf210000000000017721000000000000012000;                                                                          // add
      code[ 988] = 'h0000002400000000000001be00001500000001bd017816000000000001bf2100;                                                                          // moveLong
      code[ 989] = 'h00000023000000000000000001c02100000001a9000015000000000000000000;                                                                          // mov
      code[ 990] = 'h00000000000000000000000001c121000000000001c021000000000000012000;                                                                          // add
      code[ 991] = 'h00000023000000000000000001c22100000001a9000615000000000000000000;                                                                          // mov
      code[ 992] = 'h0000002000000000000000000000010000000000007520000000000000000000;                                                                          // label
      code[ 993] = 'h00000023000000000000000001c3210000000000000020000000000000000000;                                                                          // mov
      code[ 994] = 'h0000002000000000000000000000010000000000007620000000000000000000;                                                                          // label
      code[ 995] = 'h000000190000000000000006007821000000000001c321000000000001c12100;                                                                          // jGe
      code[ 996] = 'h00000023000000000000000001c42100000001c201c316000000000000000000;                                                                          // mov
      code[ 997] = 'h0000002300000000000001c4000215000000000001a921000000000000000000;                                                                          // mov
      code[ 998] = 'h0000002000000000000000000000010000000000007720000000000000000000;                                                                          // label
      code[ 999] = 'h00000000000000000000000001c321000000000001c321000000000000012000;                                                                          // add
      code[1000] = 'h0000001f00000000fffffffa0076210000000000000000000000000000000000;                                                                          // jmp
      code[1001] = 'h0000002000000000000000000000010000000000007820000000000000000000;                                                                          // label
      code[1002] = 'h00000023000000000000000001c52100000001ac000015000000000000000000;                                                                          // mov
      code[1003] = 'h00000000000000000000000001c621000000000001c521000000000000012000;                                                                          // add
      code[1004] = 'h00000023000000000000000001c72100000001ac000615000000000000000000;                                                                          // mov
      code[1005] = 'h0000002000000000000000000000010000000000007920000000000000000000;                                                                          // label
      code[1006] = 'h00000023000000000000000001c8210000000000000020000000000000000000;                                                                          // mov
      code[1007] = 'h0000002000000000000000000000010000000000007a20000000000000000000;                                                                          // label
      code[1008] = 'h000000190000000000000006007c21000000000001c821000000000001c62100;                                                                          // jGe
      code[1009] = 'h00000023000000000000000001c92100000001c701c816000000000000000000;                                                                          // mov
      code[1010] = 'h0000002300000000000001c9000215000000000001ac21000000000000000000;                                                                          // mov
      code[1011] = 'h0000002000000000000000000000010000000000007b20000000000000000000;                                                                          // label
      code[1012] = 'h00000000000000000000000001c821000000000001c821000000000000012000;                                                                          // add
      code[1013] = 'h0000001f00000000fffffffa007a210000000000000000000000000000000000;                                                                          // jmp
      code[1014] = 'h0000002000000000000000000000010000000000007c20000000000000000000;                                                                          // label
      code[1015] = 'h0000001f00000000000000100074210000000000000000000000000000000000;                                                                          // jmp
      code[1016] = 'h0000002000000000000000000000010000000000007320000000000000000000;                                                                          // label
      code[1017] = 'h00000001000000000000000001ca210000000000000820000000000000000000;                                                                          // array
      code[1018] = 'h00000023000000000000016a000615000000000001ca21000000000000000000;                                                                          // mov
      code[1019] = 'h00000023000000000000000001cb21000000016a000415000000000000000000;                                                                          // mov
      code[1020] = 'h00000023000000000000000001cc2100000001a9000415000000000000000000;                                                                          // mov
      code[1021] = 'h0000002400000000000001cc00001500000001cb000015000000000001772100;                                                                          // moveLong
      code[1022] = 'h00000023000000000000000001cd21000000016a000515000000000000000000;                                                                          // mov
      code[1023] = 'h00000023000000000000000001ce2100000001a9000515000000000000000000;                                                                          // mov
      code[1024] = 'h0000002400000000000001ce00001500000001cd000015000000000001772100;                                                                          // moveLong
      code[1025] = 'h00000023000000000000000001cf21000000016a000415000000000000000000;                                                                          // mov
      code[1026] = 'h00000023000000000000000001d02100000001ac000415000000000000000000;                                                                          // mov
      code[1027] = 'h0000002400000000000001d000001500000001cf017816000000000001772100;                                                                          // moveLong
      code[1028] = 'h00000023000000000000000001d121000000016a000515000000000000000000;                                                                          // mov
      code[1029] = 'h00000023000000000000000001d22100000001ac000515000000000000000000;                                                                          // mov
      code[1030] = 'h0000002400000000000001d200001500000001d1017816000000000001772100;                                                                          // moveLong
      code[1031] = 'h0000002000000000000000000000010000000000007420000000000000000000;                                                                          // label
      code[1032] = 'h0000002300000000000001a90002150000000000016a21000000000000000000;                                                                          // mov
      code[1033] = 'h0000002300000000000001ac0002150000000000016a21000000000000000000;                                                                          // mov
      code[1034] = 'h00000023000000000000000001d321000000016a000415000000000000000000;                                                                          // mov
      code[1035] = 'h00000023000000000000000001d42100000001d3017716000000000000000000;                                                                          // mov
      code[1036] = 'h00000023000000000000000001d521000000016a000515000000000000000000;                                                                          // mov
      code[1037] = 'h00000023000000000000000001d62100000001d5017716000000000000000000;                                                                          // mov
      code[1038] = 'h00000023000000000000000001d721000000016a000415000000000000000000;                                                                          // mov
      code[1039] = 'h0000002300000000000001d7000015000000000001d421000000000000000000;                                                                          // mov
      code[1040] = 'h00000023000000000000000001d821000000016a000515000000000000000000;                                                                          // mov
      code[1041] = 'h0000002300000000000001d8000015000000000001d621000000000000000000;                                                                          // mov
      code[1042] = 'h00000023000000000000000001d921000000016a000615000000000000000000;                                                                          // mov
      code[1043] = 'h0000002300000000000001d9000015000000000001a921000000000000000000;                                                                          // mov
      code[1044] = 'h00000023000000000000000001da21000000016a000615000000000000000000;                                                                          // mov
      code[1045] = 'h0000002300000000000001da000115000000000001ac21000000000000000000;                                                                          // mov
      code[1046] = 'h00000023000000000000016a0000150000000000000120000000000000000000;                                                                          // mov
      code[1047] = 'h00000023000000000000000001db21000000016a000415000000000000000000;                                                                          // mov
      code[1048] = 'h00000031000000000000000001db210000000000000120000000000000062000;                                                                          // resize
      code[1049] = 'h00000023000000000000000001dc21000000016a000515000000000000000000;                                                                          // mov
      code[1050] = 'h00000031000000000000000001dc210000000000000120000000000000072000;                                                                          // resize
      code[1051] = 'h00000023000000000000000001dd21000000016a000615000000000000000000;                                                                          // mov
      code[1052] = 'h00000031000000000000000001dd210000000000000220000000000000082000;                                                                          // resize
      code[1053] = 'h0000001f00000000000000020067210000000000000000000000000000000000;                                                                          // jmp
      code[1054] = 'h0000001f00000000000000060069210000000000000000000000000000000000;                                                                          // jmp
      code[1055] = 'h0000002000000000000000000000010000000000006720000000000000000000;                                                                          // label
      code[1056] = 'h0000002300000000000000000173210000000000000120000000000000000000;                                                                          // mov
      code[1057] = 'h0000001f00000000000000030069210000000000000000000000000000000000;                                                                          // jmp
      code[1058] = 'h0000002000000000000000000000010000000000006820000000000000000000;                                                                          // label
      code[1059] = 'h0000002300000000000000000173210000000000000020000000000000000000;                                                                          // mov
      code[1060] = 'h0000002000000000000000000000010000000000006920000000000000000000;                                                                          // label
      code[1061] = 'h0000002000000000000000000000010000000000000720000000000000000000;                                                                          // label
      code[1062] = 'h0000002000000000000000000000010000000000000820000000000000000000;                                                                          // label
      code[1063] = 'h0000002000000000000000000000010000000000000920000000000000000000;                                                                          // label
      code[1064] = 'h0000001400000000000000000006210000000000000320000000000000000000;                                                                          // free
      code[1065] = 'h0000001f00000000000000490002210000000000000000000000000000000000;                                                                          // jmp
      code[1066] = 'h0000002000000000000000000000010000000000000520000000000000000000;                                                                          // label
      code[1067] = 'h0000001d0000000000000045007d210000000000000221000000000000022000;                                                                          // jNe
      code[1068] = 'h00000015000000000000000001de210000000000000000000000000000000000;                                                                          // in
      code[1069] = 'h0000002000000000000000000000010000000000007e20000000000000000000;                                                                          // label
      code[1070] = 'h00000023000000000000000001df210000000003000315000000000000000000;                                                                          // mov
      code[1071] = 'h0000001d0000000000000005008221000000000001df21000000000000002000;                                                                          // jNe
      code[1072] = 'h000000230000000000000000000015000000000001df21000000000000000000;                                                                          // mov
      code[1073] = 'h0000002300000000000000000001150000000000000320000000000000000000;                                                                          // mov
      code[1074] = 'h0000002300000000000000000002150000000000000020000000000000000000;                                                                          // mov
      code[1075] = 'h0000001f000000000000002f0081210000000000000000000000000000000000;                                                                          // jmp
      code[1076] = 'h0000002000000000000000000000010000000000008220000000000000000000;                                                                          // label
      code[1077] = 'h0000002000000000000000000000010000000000008320000000000000000000;                                                                          // label
      code[1078] = 'h00000023000000000000000001e0210000000000000020000000000000000000;                                                                          // mov
      code[1079] = 'h0000002000000000000000000000010000000000008420000000000000000000;                                                                          // label
      code[1080] = 'h000000190000000000000026008621000000000001e021000000000000632000;                                                                          // jGe
      code[1081] = 'h00000039000000000000000001e12100000001df000015000000000000012000;                                                                          // subtract
      code[1082] = 'h00000023000000000000000001e22100000001df000415000000000000000000;                                                                          // mov
      code[1083] = 'h0000001b000000000000000d008721000000000001de2100000001e201e11600;                                                                          // jLe
      code[1084] = 'h00000000000000000000000001e321000000000001e121000000000000012000;                                                                          // add
      code[1085] = 'h00000026000000000000000001e42100000001df000615000000000000000000;                                                                          // not
      code[1086] = 'h000000170000000000000005008821000000000001e421000000000000002000;                                                                          // jEq
      code[1087] = 'h000000230000000000000000000015000000000001df21000000000000000000;                                                                          // mov
      code[1088] = 'h0000002300000000000000000001150000000000000220000000000000000000;                                                                          // mov
      code[1089] = 'h000000230000000000000000000215000000000001e321000000000000000000;                                                                          // mov
      code[1090] = 'h0000001f00000000000000200081210000000000000000000000000000000000;                                                                          // jmp
      code[1091] = 'h0000002000000000000000000000010000000000008820000000000000000000;                                                                          // label
      code[1092] = 'h00000023000000000000000001e52100000001df000615000000000000000000;                                                                          // mov
      code[1093] = 'h00000023000000000000000001e62100000001e501e316000000000000000000;                                                                          // mov
      code[1094] = 'h00000023000000000000000001df21000000000001e621000000000000000000;                                                                          // mov
      code[1095] = 'h0000001f00000000000000140085210000000000000000000000000000000000;                                                                          // jmp
      code[1096] = 'h0000002000000000000000000000010000000000008720000000000000000000;                                                                          // label
      code[1097] = 'h00000005000000000000000001e721000000000001e221000000000001de2100;                                                                          // arrayIndex
      code[1098] = 'h000000170000000000000005008921000000000001e721000000000000002000;                                                                          // jEq
      code[1099] = 'h000000230000000000000000000015000000000001df21000000000000000000;                                                                          // mov
      code[1100] = 'h0000002300000000000000000001150000000000000120000000000000000000;                                                                          // mov
      code[1101] = 'h000000390000000000000000000215000000000001e721000000000000012000;                                                                          // subtract
      code[1102] = 'h0000001f00000000000000140081210000000000000000000000000000000000;                                                                          // jmp
      code[1103] = 'h0000002000000000000000000000010000000000008920000000000000000000;                                                                          // label
      code[1104] = 'h00000003000000000000000001e821000000000001e221000000000001de2100;                                                                          // arrayCountLess
      code[1105] = 'h00000026000000000000000001e92100000001df000615000000000000000000;                                                                          // not
      code[1106] = 'h000000170000000000000005008a21000000000001e921000000000000002000;                                                                          // jEq
      code[1107] = 'h000000230000000000000000000015000000000001df21000000000000000000;                                                                          // mov
      code[1108] = 'h0000002300000000000000000001150000000000000020000000000000000000;                                                                          // mov
      code[1109] = 'h000000230000000000000000000215000000000001e821000000000000000000;                                                                          // mov
      code[1110] = 'h0000001f000000000000000c0081210000000000000000000000000000000000;                                                                          // jmp
      code[1111] = 'h0000002000000000000000000000010000000000008a20000000000000000000;                                                                          // label
      code[1112] = 'h00000023000000000000000001ea2100000001df000615000000000000000000;                                                                          // mov
      code[1113] = 'h00000023000000000000000001eb2100000001ea01e816000000000000000000;                                                                          // mov
      code[1114] = 'h00000023000000000000000001df21000000000001eb21000000000000000000;                                                                          // mov
      code[1115] = 'h0000002000000000000000000000010000000000008520000000000000000000;                                                                          // label
      code[1116] = 'h00000000000000000000000001e021000000000001e021000000000000012000;                                                                          // add
      code[1117] = 'h0000001f00000000ffffffda0084210000000000000000000000000000000000;                                                                          // jmp
      code[1118] = 'h0000002000000000000000000000010000000000008620000000000000000000;                                                                          // label
      code[1119] = 'h0000000800000000000000000000010000000000000000000000000000000000;                                                                          // assert
      code[1120] = 'h0000002000000000000000000000010000000000007f20000000000000000000;                                                                          // label
      code[1121] = 'h0000002000000000000000000000010000000000008020000000000000000000;                                                                          // label
      code[1122] = 'h0000002000000000000000000000010000000000008120000000000000000000;                                                                          // label
      code[1123] = 'h00000023000000000000000001ec210000000000000115000000000000000000;                                                                          // mov
      code[1124] = 'h0000001d0000000000000008008b21000000000001ec21000000000000012000;                                                                          // jNe
      code[1125] = 'h0000002700000000000000000000010000000000000120000000000000000000;                                                                          // out
      code[1126] = 'h00000023000000000000000001ed210000000000000015000000000000000000;                                                                          // mov
      code[1127] = 'h00000023000000000000000001ee210000000000000215000000000000000000;                                                                          // mov
      code[1128] = 'h00000023000000000000000001ef2100000001ed000515000000000000000000;                                                                          // mov
      code[1129] = 'h00000023000000000000000001f02100000001ef01ee16000000000000000000;                                                                          // mov
      code[1130] = 'h000000270000000000000000000001000000000001f021000000000000000000;                                                                          // out
      code[1131] = 'h0000001f0000000000000003008c210000000000000000000000000000000000;                                                                          // jmp
      code[1132] = 'h0000002000000000000000000000010000000000008b20000000000000000000;                                                                          // label
      code[1133] = 'h0000002700000000000000000000010000000000000020000000000000000000;                                                                          // out
      code[1134] = 'h0000002000000000000000000000010000000000008c20000000000000000000;                                                                          // label
      code[1135] = 'h0000001f00000000000000030002210000000000000000000000000000000000;                                                                          // jmp
      code[1136] = 'h0000002000000000000000000000010000000000007d20000000000000000000;                                                                          // label
      code[1137] = 'h0000001f00000000000000030003210000000000000000000000000000000000;                                                                          // jmp
      code[1138] = 'h0000002000000000000000000000010000000000000220000000000000000000;                                                                          // label
      code[1139] = 'h0000001f00000000fffffb8e0001210000000000000000000000000000000000;                                                                          // jmp
      code[1140] = 'h0000002000000000000000000000010000000000000320000000000000000000;                                                                          // label
    end
  endtask

  task endTest();                                                               // BTree: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 0;
      success = success && outMem[1] == 1;
      success = success && outMem[2] == 22;
      success = success && outMem[3] == 0;
      success = success && outMem[4] == 1;
      success = success && outMem[5] == 33;
    end
  endtask
