  parameter integer NInstructions = 6;

  task startTest();                                                             // Not_test: load code
    begin

      code[   0] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   1] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[   2] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000001000000100001000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[   3] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   4] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   5] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
    end
  endtask

  task endTest();                                                               // Not_test: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 3;
      success = success && outMem[1] == 0;
      success = success && outMem[2] == 1;
    end
  endtask
