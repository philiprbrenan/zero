  parameter integer NInstructions = 7;

  task startTest();                                                             // Pop_test: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000110000000000010000000000;                                          // push
      code[   2] = 'b0000000000000000000000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000110000000000010000000000;                                          // push
      code[   3] = 'b0000000000000000000000001011010000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000110000000000010000000000;                                          // pop
      code[   4] = 'b0000000000000000000000001011010000000000000000000000000000000000000000000000000000000000000000000000000001000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000110000000000010000000000;                                          // pop
      code[   5] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   6] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
    end
  endtask

  task endTest();                                                               // Pop_test: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 2;
      success = success && outMem[1] == 1;
    end
  endtask
