  parameter integer NInstructions = 28;

  task startTest();                                                             // Array_scans: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   2] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000000010100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   3] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000000000000111100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   4] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000011110000000010000000000;                                          // arrayIndex
      code[   5] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   6] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000001000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000001010000000010000000000;                                          // arrayIndex
      code[   7] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   8] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000011000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000010100000000010000000000;                                          // arrayIndex
      code[   9] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  10] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000100000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000111100000000010000000000;                                          // arrayIndex
      code[  11] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  12] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000010100000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000110001000000010000000000;                                          // arrayCountLess
      code[  13] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  14] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000001100000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000100110000000010000000000;                                          // arrayCountLess
      code[  15] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  16] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000011100000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000111100000000010000000000;                                          // arrayCountLess
      code[  17] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  18] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000010000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000101000000000010000000000;                                          // arrayCountLess
      code[  19] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  20] = 'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010010000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000110001000000010000000000;                                          // arrayCountGreater
      code[  21] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  22] = 'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001010000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000100110000000010000000000;                                          // arrayCountGreater
      code[  23] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  24] = 'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000011010000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000111100000000010000000000;                                          // arrayCountGreater
      code[  25] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  26] = 'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000110000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000101000000000010000000000;                                          // arrayCountGreater
      code[  27] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
    end
  endtask

  task endTest();                                                               // Array_scans: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 3;
      success = success && outMem[1] == 2;
      success = success && outMem[2] == 1;
      success = success && outMem[3] == 0;
      success = success && outMem[4] == 3;
      success = success && outMem[5] == 2;
      success = success && outMem[6] == 1;
      success = success && outMem[7] == 0;
      success = success && outMem[8] == 0;
      success = success && outMem[9] == 1;
      success = success && outMem[10] == 2;
      success = success && outMem[11] == 3;
    end
  endtask
