  task startTest();                                                             // Jeq_test: load code
    begin
      NInstructionEnd = 12;

      code[   0] = 'h0000002000000000000000000000010000000000000120000000000000000000;                                                                          // label
      code[   1] = 'h0000002300000000000000000000210000000000000120000000000000000000;                                                                          // mov
      code[   2] = 'h0000002300000000000000000001210000000000000220000000000000000000;                                                                          // mov
      code[   3] = 'h0000001700000000000000050002210000000000000021000000000000012100;                                                                          // jEq
      code[   4] = 'h0000002700000000000000000000010000000000006f20000000000000000000;                                                                          // out
      code[   5] = 'h0000001700000000000000030002210000000000000021000000000000002100;                                                                          // jEq
      code[   6] = 'h000000270000000000000000000001000000000000de20000000000000000000;                                                                          // out
      code[   7] = 'h0000001f00000000000000040004210000000000000000000000000000000000;                                                                          // jmp
      code[   8] = 'h0000002000000000000000000000010000000000000220000000000000000000;                                                                          // label
      code[   9] = 'h0000002700000000000000000000010000000000014d20000000000000000000;                                                                          // out
      code[  10] = 'h0000002000000000000000000000010000000000000320000000000000000000;                                                                          // label
      code[  11] = 'h0000002000000000000000000000010000000000000420000000000000000000;                                                                          // label
    end
  endtask

  task endTest();                                                               // Jeq_test: Evaluate results in out channel
    begin
      success = 1;

    end
  endtask
