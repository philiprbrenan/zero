  parameter integer NInstructions = 5;

  task startTest();                                                             // Shift_up_test: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   2] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   3] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   4] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000001100011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
    end
  endtask

  task endTest();                                                               // Shift_up_test: Evaluate results in out channel
    begin
      success = 1;
    end
  endtask
