//-----------------------------------------------------------------------------
// Fpga test
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
module fpga                                                                     // Run test programs
 (input  wire run,                                                              // Run - clock at lest once to allow code to be loaded
  output reg  finished,                                                         // Goes high when the program has finished
  output reg  success);                                                         // Goes high on finish if all the tests passed

  parameter integer MemoryElementWidth =  12;                                   // Memory element width

  parameter integer NArea   =        7;                                         // Size of each area on the heap
  parameter integer NArrays =       15;                                         // Maximum number of arrays
  parameter integer NHeap   =      105;                                         // Amount of heap memory
  parameter integer NLocal  =     2748;                                         // Size of local memory
  parameter integer NOut    =        0;                                         // Size of output area
  parameter integer NIn     =        0;                                         // Size of input area
  reg [MemoryElementWidth-1:0]   arraySizes[NArrays-1:0];                       // Size of each array
  reg [MemoryElementWidth-1:0]      heapMem[NHeap-1  :0];                       // Heap memory
  reg [MemoryElementWidth-1:0]     localMem[NLocal-1 :0];                       // Local memory
  reg [MemoryElementWidth-1:0]       outMem[NOut-1   :0];                       // Out channel
  reg [MemoryElementWidth-1:0]        inMem[NIn-1    :0];                       // In channel
  reg [MemoryElementWidth-1:0]  freedArrays[NArrays-1:0];                       // Freed arrays list implemented as a stack
  reg [MemoryElementWidth-1:0]   arrayShift[NArea-1  :0];                       // Array shift area

  integer inMemPos;                                                             // Current position in input channel
  integer outMemPos;                                                            // Position in output channel
  integer allocs;                                                               // Maximum number of array allocations in use at any one time
  integer freedArraysTop;                                                       // Position in freed arrays stack

  integer ip;                                                                   // Instruction pointer
  reg     clock;                                                                // Clock - has to be one bit wide for yosys
  integer steps;                                                                // Number of steps executed so far
  integer i, j, k;                                                              // A useful counter

  task updateArrayLength(input integer arena, input integer array, input integer index); // Update array length if we are updating an array
    begin
      if (arena == 1 && arraySizes[array] < index + 1) arraySizes[array] = index + 1;
    end
  endtask

  always @(posedge run) begin                                                   // Initialize
    ip             = 0;
    clock          = 0;
    steps          = 0;
    finished       = 0;
    success        = 0;
    inMemPos       = 0;
    outMemPos      = 0;
    allocs         = 0;
    freedArraysTop = 0;
    if (0) begin                                                  // Clear memory
      for(i = 0; i < NHeap;   i = i + 1)    heapMem[i] = 0;
      for(i = 0; i < NLocal;  i = i + 1)   localMem[i] = 0;
      for(i = 0; i < NArrays; i = i + 1) arraySizes[i] = 0;
    end
  end

  always @(clock) begin                                                         // Each instruction
    steps = steps + 1;
    case(ip)

          0 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[0] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[0] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[0]] = 0;
              ip = 1;
      end

          1 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*7 + 2] = 3;
              updateArrayLength(1, localMem[0], 2);
              ip = 2;
      end

          2 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*7 + 3] = 0;
              updateArrayLength(1, localMem[0], 3);
              ip = 3;
      end

          3 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = 0;
              updateArrayLength(1, localMem[0], 0);
              ip = 4;
      end

          4 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*7 + 1] = 0;
              updateArrayLength(1, localMem[0], 1);
              ip = 5;
      end

          5 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1]] = 0;
              ip = 6;
      end

          6 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 7;
      end

          7 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 8;
      end

          8 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2] != 0 ? 31 : 9;
      end

          9 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[3] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[3] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[3]] = 0;
              ip = 10;
      end

         10 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 0] = 1;
              updateArrayLength(1, localMem[3], 0);
              ip = 11;
      end

         11 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 2] = 0;
              updateArrayLength(1, localMem[3], 2);
              ip = 12;
      end

         12 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[4] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[4] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[4]] = 0;
              ip = 13;
      end

         13 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 4] = localMem[4];
              updateArrayLength(1, localMem[3], 4);
              ip = 14;
      end

         14 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[5] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[5] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[5]] = 0;
              ip = 15;
      end

         15 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 5] = localMem[5];
              updateArrayLength(1, localMem[3], 5);
              ip = 16;
      end

         16 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 6] = 0;
              updateArrayLength(1, localMem[3], 6);
              ip = 17;
      end

         17 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 3] = localMem[0];
              updateArrayLength(1, localMem[3], 3);
              ip = 18;
      end

         18 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 1] = heapMem[localMem[0]*7 + 1] + 1;
              updateArrayLength(1, localMem[0], 1);
              ip = 19;
      end

         19 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[3]*7 + 1] = heapMem[localMem[0]*7 + 1];
              updateArrayLength(1, localMem[3], 1);
              ip = 20;
      end

         20 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[6] = heapMem[localMem[3]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 21;
      end

         21 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[6]*7 + 0] = 1;
              updateArrayLength(1, localMem[6], 0);
              ip = 22;
      end

         22 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[7] = heapMem[localMem[3]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 23;
      end

         23 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[7]*7 + 0] = 11;
              updateArrayLength(1, localMem[7], 0);
              ip = 24;
      end

         24 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = heapMem[localMem[0]*7 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 25;
      end

         25 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[0]*7 + 3] = localMem[3];
              updateArrayLength(1, localMem[0], 3);
              ip = 26;
      end

         26 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[8] = heapMem[localMem[3]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 27;
      end

         27 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[8]] = 1;
              ip = 28;
      end

         28 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[9] = heapMem[localMem[3]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 29;
      end

         29 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[9]] = 1;
              ip = 30;
      end

         30 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 1059;
      end

         31 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    31");
      end

         32 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    32");
      end

         33 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    33");
      end

         34 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed    34");
      end

         35 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    35");
      end

         36 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed    36");
      end

         37 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed    37");
      end

         38 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed    38");
      end

         39 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    39");
      end

         40 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed    40");
      end

         41 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed    41");
      end

         42 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed    42");
      end

         43 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    43");
      end

         44 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    44");
      end

         45 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed    45");
      end

         46 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    46");
      end

         47 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed    47");
      end

         48 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    48");
      end

         49 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed    49");
      end

         50 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
         $display("Should not be executed    50");
      end

         51 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed    51");
      end

         52 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    52");
      end

         53 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    53");
      end

         54 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    54");
      end

         55 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    55");
      end

         56 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed    56");
      end

         57 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed    57");
      end

         58 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed    58");
      end

         59 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    59");
      end

         60 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed    60");
      end

         61 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    61");
      end

         62 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed    62");
      end

         63 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    63");
      end

         64 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed    64");
      end

         65 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed    65");
      end

         66 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed    66");
      end

         67 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed    67");
      end

         68 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    68");
      end

         69 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    69");
      end

         70 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    70");
      end

         71 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    71");
      end

         72 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed    72");
      end

         73 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    73");
      end

         74 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    74");
      end

         75 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    75");
      end

         76 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed    76");
      end

         77 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    77");
      end

         78 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed    78");
      end

         79 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed    79");
      end

         80 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    80");
      end

         81 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed    81");
      end

         82 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed    82");
      end

         83 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    83");
      end

         84 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    84");
      end

         85 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed    85");
      end

         86 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    86");
      end

         87 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed    87");
      end

         88 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    88");
      end

         89 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    89");
      end

         90 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    90");
      end

         91 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed    91");
      end

         92 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    92");
      end

         93 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed    93");
      end

         94 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed    94");
      end

         95 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed    95");
      end

         96 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    96");
      end

         97 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    97");
      end

         98 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed    98");
      end

         99 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed    99");
      end

        100 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   100");
      end

        101 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   101");
      end

        102 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   102");
      end

        103 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   103");
      end

        104 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   104");
      end

        105 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   105");
      end

        106 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   106");
      end

        107 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   107");
      end

        108 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   108");
      end

        109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   109");
      end

        110 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   110");
      end

        111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   111");
      end

        112 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   112");
      end

        113 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   113");
      end

        114 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   114");
      end

        115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   115");
      end

        116 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   116");
      end

        117 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   117");
      end

        118 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   118");
      end

        119 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   119");
      end

        120 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   120");
      end

        121 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   121");
      end

        122 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   122");
      end

        123 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   123");
      end

        124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   124");
      end

        125 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   125");
      end

        126 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   126");
      end

        127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   127");
      end

        128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   128");
      end

        129 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   129");
      end

        130 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   130");
      end

        131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   131");
      end

        132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   132");
      end

        133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   133");
      end

        134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   134");
      end

        135 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   135");
      end

        136 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   136");
      end

        137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   137");
      end

        138 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   138");
      end

        139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   139");
      end

        140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   140");
      end

        141 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   141");
      end

        142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   142");
      end

        143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   143");
      end

        144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   144");
      end

        145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   145");
      end

        146 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   146");
      end

        147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   147");
      end

        148 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   148");
      end

        149 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   149");
      end

        150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   150");
      end

        151 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   151");
      end

        152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   152");
      end

        153 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   153");
      end

        154 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   154");
      end

        155 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   155");
      end

        156 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed   156");
      end

        157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   157");
      end

        158 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed   158");
      end

        159 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   159");
      end

        160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   160");
      end

        161 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   161");
      end

        162 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   162");
      end

        163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   163");
      end

        164 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   164");
      end

        165 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   165");
      end

        166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   166");
      end

        167 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   167");
      end

        168 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   168");
      end

        169 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   169");
      end

        170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   170");
      end

        171 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   171");
      end

        172 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   172");
      end

        173 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   173");
      end

        174 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   174");
      end

        175 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   175");
      end

        176 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   176");
      end

        177 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   177");
      end

        178 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   178");
      end

        179 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   179");
      end

        180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   180");
      end

        181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   181");
      end

        182 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   182");
      end

        183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   183");
      end

        184 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   184");
      end

        185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   185");
      end

        186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   186");
      end

        187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   187");
      end

        188 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   188");
      end

        189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   189");
      end

        190 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   190");
      end

        191 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   191");
      end

        192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   192");
      end

        193 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   193");
      end

        194 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   194");
      end

        195 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   195");
      end

        196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   196");
      end

        197 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   197");
      end

        198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   198");
      end

        199 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   199");
      end

        200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   200");
      end

        201 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   201");
      end

        202 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   202");
      end

        203 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   203");
      end

        204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   204");
      end

        205 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   205");
      end

        206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   206");
      end

        207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   207");
      end

        208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   208");
      end

        209 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   209");
      end

        210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   210");
      end

        211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   211");
      end

        212 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   212");
      end

        213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   213");
      end

        214 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   214");
      end

        215 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   215");
      end

        216 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   216");
      end

        217 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   217");
      end

        218 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   218");
      end

        219 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   219");
      end

        220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   220");
      end

        221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   221");
      end

        222 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   222");
      end

        223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   223");
      end

        224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   224");
      end

        225 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   225");
      end

        226 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   226");
      end

        227 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   227");
      end

        228 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   228");
      end

        229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   229");
      end

        230 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   230");
      end

        231 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   231");
      end

        232 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   232");
      end

        233 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   233");
      end

        234 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   234");
      end

        235 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   235");
      end

        236 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   236");
      end

        237 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   237");
      end

        238 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   238");
      end

        239 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   239");
      end

        240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   240");
      end

        241 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   241");
      end

        242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   242");
      end

        243 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   243");
      end

        244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   244");
      end

        245 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   245");
      end

        246 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   246");
      end

        247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   247");
      end

        248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   248");
      end

        249 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   249");
      end

        250 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   250");
      end

        251 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   251");
      end

        252 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   252");
      end

        253 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   253");
      end

        254 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   254");
      end

        255 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   255");
      end

        256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   256");
      end

        257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   257");
      end

        258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   258");
      end

        259 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   259");
      end

        260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   260");
      end

        261 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   261");
      end

        262 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   262");
      end

        263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   263");
      end

        264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   264");
      end

        265 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   265");
      end

        266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   266");
      end

        267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   267");
      end

        268 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   268");
      end

        269 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   269");
      end

        270 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   270");
      end

        271 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   271");
      end

        272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   272");
      end

        273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   273");
      end

        274 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   274");
      end

        275 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   275");
      end

        276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   276");
      end

        277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   277");
      end

        278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   278");
      end

        279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   279");
      end

        280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   280");
      end

        281 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   281");
      end

        282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   282");
      end

        283 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   283");
      end

        284 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   284");
      end

        285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   285");
      end

        286 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   286");
      end

        287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   287");
      end

        288 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   288");
      end

        289 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   289");
      end

        290 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   290");
      end

        291 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   291");
      end

        292 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   292");
      end

        293 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   293");
      end

        294 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   294");
      end

        295 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   295");
      end

        296 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   296");
      end

        297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   297");
      end

        298 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   298");
      end

        299 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   299");
      end

        300 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   300");
      end

        301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   301");
      end

        302 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   302");
      end

        303 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   303");
      end

        304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   304");
      end

        305 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   305");
      end

        306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   306");
      end

        307 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   307");
      end

        308 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
         $display("Should not be executed   308");
      end

        309 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   309");
      end

        310 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed   310");
      end

        311 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   311");
      end

        312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   312");
      end

        313 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   313");
      end

        314 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   314");
      end

        315 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   315");
      end

        316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   316");
      end

        317 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   317");
      end

        318 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   318");
      end

        319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   319");
      end

        320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   320");
      end

        321 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   321");
      end

        322 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed   322");
      end

        323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   323");
      end

        324 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed   324");
      end

        325 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   325");
      end

        326 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   326");
      end

        327 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed   327");
      end

        328 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   328");
      end

        329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   329");
      end

        330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   330");
      end

        331 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   331");
      end

        332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   332");
      end

        333 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   333");
      end

        334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   334");
      end

        335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   335");
      end

        336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   336");
      end

        337 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   337");
      end

        338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   338");
      end

        339 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   339");
      end

        340 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   340");
      end

        341 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   341");
      end

        342 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   342");
      end

        343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   343");
      end

        344 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   344");
      end

        345 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   345");
      end

        346 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   346");
      end

        347 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   347");
      end

        348 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   348");
      end

        349 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   349");
      end

        350 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   350");
      end

        351 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   351");
      end

        352 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   352");
      end

        353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   353");
      end

        354 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   354");
      end

        355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   355");
      end

        356 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   356");
      end

        357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   357");
      end

        358 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   358");
      end

        359 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   359");
      end

        360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   360");
      end

        361 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   361");
      end

        362 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   362");
      end

        363 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   363");
      end

        364 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   364");
      end

        365 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   365");
      end

        366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   366");
      end

        367 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   367");
      end

        368 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   368");
      end

        369 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   369");
      end

        370 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   370");
      end

        371 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   371");
      end

        372 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   372");
      end

        373 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   373");
      end

        374 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   374");
      end

        375 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   375");
      end

        376 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   376");
      end

        377 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   377");
      end

        378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   378");
      end

        379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   379");
      end

        380 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   380");
      end

        381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   381");
      end

        382 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   382");
      end

        383 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   383");
      end

        384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   384");
      end

        385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   385");
      end

        386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   386");
      end

        387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   387");
      end

        388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   388");
      end

        389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   389");
      end

        390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   390");
      end

        391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   391");
      end

        392 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   392");
      end

        393 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   393");
      end

        394 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   394");
      end

        395 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   395");
      end

        396 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   396");
      end

        397 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   397");
      end

        398 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   398");
      end

        399 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   399");
      end

        400 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   400");
      end

        401 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   401");
      end

        402 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed   402");
      end

        403 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   403");
      end

        404 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed   404");
      end

        405 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   405");
      end

        406 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   406");
      end

        407 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   407");
      end

        408 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   408");
      end

        409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   409");
      end

        410 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   410");
      end

        411 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   411");
      end

        412 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   412");
      end

        413 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   413");
      end

        414 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   414");
      end

        415 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   415");
      end

        416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   416");
      end

        417 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   417");
      end

        418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   418");
      end

        419 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   419");
      end

        420 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   420");
      end

        421 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   421");
      end

        422 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   422");
      end

        423 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   423");
      end

        424 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   424");
      end

        425 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   425");
      end

        426 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   426");
      end

        427 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   427");
      end

        428 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   428");
      end

        429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   429");
      end

        430 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   430");
      end

        431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   431");
      end

        432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   432");
      end

        433 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   433");
      end

        434 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   434");
      end

        435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   435");
      end

        436 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   436");
      end

        437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   437");
      end

        438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   438");
      end

        439 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   439");
      end

        440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   440");
      end

        441 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   441");
      end

        442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   442");
      end

        443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   443");
      end

        444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   444");
      end

        445 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   445");
      end

        446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   446");
      end

        447 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   447");
      end

        448 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   448");
      end

        449 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   449");
      end

        450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   450");
      end

        451 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   451");
      end

        452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   452");
      end

        453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   453");
      end

        454 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   454");
      end

        455 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   455");
      end

        456 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   456");
      end

        457 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   457");
      end

        458 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   458");
      end

        459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   459");
      end

        460 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   460");
      end

        461 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   461");
      end

        462 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   462");
      end

        463 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   463");
      end

        464 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   464");
      end

        465 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   465");
      end

        466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   466");
      end

        467 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   467");
      end

        468 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   468");
      end

        469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   469");
      end

        470 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   470");
      end

        471 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   471");
      end

        472 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   472");
      end

        473 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   473");
      end

        474 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   474");
      end

        475 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   475");
      end

        476 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   476");
      end

        477 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   477");
      end

        478 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   478");
      end

        479 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   479");
      end

        480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   480");
      end

        481 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   481");
      end

        482 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   482");
      end

        483 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   483");
      end

        484 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   484");
      end

        485 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   485");
      end

        486 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   486");
      end

        487 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   487");
      end

        488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   488");
      end

        489 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   489");
      end

        490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   490");
      end

        491 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   491");
      end

        492 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   492");
      end

        493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   493");
      end

        494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   494");
      end

        495 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   495");
      end

        496 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   496");
      end

        497 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   497");
      end

        498 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   498");
      end

        499 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   499");
      end

        500 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   500");
      end

        501 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   501");
      end

        502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   502");
      end

        503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   503");
      end

        504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   504");
      end

        505 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   505");
      end

        506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   506");
      end

        507 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   507");
      end

        508 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   508");
      end

        509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   509");
      end

        510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   510");
      end

        511 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   511");
      end

        512 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   512");
      end

        513 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   513");
      end

        514 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   514");
      end

        515 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   515");
      end

        516 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   516");
      end

        517 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   517");
      end

        518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   518");
      end

        519 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   519");
      end

        520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   520");
      end

        521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   521");
      end

        522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   522");
      end

        523 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   523");
      end

        524 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   524");
      end

        525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   525");
      end

        526 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   526");
      end

        527 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   527");
      end

        528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   528");
      end

        529 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   529");
      end

        530 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   530");
      end

        531 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   531");
      end

        532 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   532");
      end

        533 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   533");
      end

        534 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   534");
      end

        535 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   535");
      end

        536 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   536");
      end

        537 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   537");
      end

        538 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   538");
      end

        539 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   539");
      end

        540 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   540");
      end

        541 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   541");
      end

        542 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   542");
      end

        543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   543");
      end

        544 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   544");
      end

        545 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   545");
      end

        546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   546");
      end

        547 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   547");
      end

        548 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   548");
      end

        549 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   549");
      end

        550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   550");
      end

        551 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed   551");
      end

        552 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed   552");
      end

        553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   553");
      end

        554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   554");
      end

        555 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   555");
      end

        556 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   556");
      end

        557 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   557");
      end

        558 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed   558");
      end

        559 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   559");
      end

        560 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed   560");
      end

        561 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   561");
      end

        562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   562");
      end

        563 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   563");
      end

        564 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   564");
      end

        565 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   565");
      end

        566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   566");
      end

        567 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   567");
      end

        568 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   568");
      end

        569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   569");
      end

        570 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   570");
      end

        571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   571");
      end

        572 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed   572");
      end

        573 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   573");
      end

        574 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed   574");
      end

        575 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   575");
      end

        576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   576");
      end

        577 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed   577");
      end

        578 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   578");
      end

        579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   579");
      end

        580 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   580");
      end

        581 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   581");
      end

        582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   582");
      end

        583 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   583");
      end

        584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   584");
      end

        585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   585");
      end

        586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   586");
      end

        587 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   587");
      end

        588 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   588");
      end

        589 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   589");
      end

        590 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   590");
      end

        591 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   591");
      end

        592 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   592");
      end

        593 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   593");
      end

        594 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   594");
      end

        595 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   595");
      end

        596 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   596");
      end

        597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   597");
      end

        598 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   598");
      end

        599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   599");
      end

        600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   600");
      end

        601 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   601");
      end

        602 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   602");
      end

        603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   603");
      end

        604 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   604");
      end

        605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   605");
      end

        606 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   606");
      end

        607 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   607");
      end

        608 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   608");
      end

        609 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   609");
      end

        610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   610");
      end

        611 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   611");
      end

        612 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   612");
      end

        613 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   613");
      end

        614 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   614");
      end

        615 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   615");
      end

        616 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   616");
      end

        617 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   617");
      end

        618 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   618");
      end

        619 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   619");
      end

        620 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   620");
      end

        621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   621");
      end

        622 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   622");
      end

        623 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   623");
      end

        624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   624");
      end

        625 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   625");
      end

        626 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   626");
      end

        627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   627");
      end

        628 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   628");
      end

        629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   629");
      end

        630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   630");
      end

        631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   631");
      end

        632 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   632");
      end

        633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   633");
      end

        634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   634");
      end

        635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   635");
      end

        636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   636");
      end

        637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   637");
      end

        638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   638");
      end

        639 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   639");
      end

        640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   640");
      end

        641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   641");
      end

        642 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   642");
      end

        643 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   643");
      end

        644 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   644");
      end

        645 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   645");
      end

        646 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   646");
      end

        647 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   647");
      end

        648 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   648");
      end

        649 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   649");
      end

        650 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   650");
      end

        651 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   651");
      end

        652 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed   652");
      end

        653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   653");
      end

        654 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed   654");
      end

        655 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   655");
      end

        656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   656");
      end

        657 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   657");
      end

        658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   658");
      end

        659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   659");
      end

        660 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   660");
      end

        661 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   661");
      end

        662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   662");
      end

        663 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   663");
      end

        664 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   664");
      end

        665 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   665");
      end

        666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   666");
      end

        667 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   667");
      end

        668 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   668");
      end

        669 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   669");
      end

        670 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   670");
      end

        671 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   671");
      end

        672 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   672");
      end

        673 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   673");
      end

        674 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   674");
      end

        675 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   675");
      end

        676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   676");
      end

        677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   677");
      end

        678 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   678");
      end

        679 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   679");
      end

        680 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   680");
      end

        681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   681");
      end

        682 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   682");
      end

        683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   683");
      end

        684 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   684");
      end

        685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   685");
      end

        686 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   686");
      end

        687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   687");
      end

        688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   688");
      end

        689 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   689");
      end

        690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   690");
      end

        691 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   691");
      end

        692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   692");
      end

        693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   693");
      end

        694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   694");
      end

        695 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   695");
      end

        696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   696");
      end

        697 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   697");
      end

        698 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   698");
      end

        699 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   699");
      end

        700 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   700");
      end

        701 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   701");
      end

        702 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   702");
      end

        703 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   703");
      end

        704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   704");
      end

        705 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   705");
      end

        706 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   706");
      end

        707 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   707");
      end

        708 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   708");
      end

        709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   709");
      end

        710 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   710");
      end

        711 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   711");
      end

        712 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   712");
      end

        713 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   713");
      end

        714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   714");
      end

        715 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   715");
      end

        716 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   716");
      end

        717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   717");
      end

        718 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   718");
      end

        719 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   719");
      end

        720 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   720");
      end

        721 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   721");
      end

        722 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   722");
      end

        723 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   723");
      end

        724 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   724");
      end

        725 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   725");
      end

        726 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   726");
      end

        727 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   727");
      end

        728 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   728");
      end

        729 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   729");
      end

        730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   730");
      end

        731 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   731");
      end

        732 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   732");
      end

        733 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   733");
      end

        734 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   734");
      end

        735 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   735");
      end

        736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   736");
      end

        737 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   737");
      end

        738 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   738");
      end

        739 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   739");
      end

        740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   740");
      end

        741 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   741");
      end

        742 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   742");
      end

        743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   743");
      end

        744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   744");
      end

        745 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   745");
      end

        746 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   746");
      end

        747 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   747");
      end

        748 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   748");
      end

        749 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   749");
      end

        750 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   750");
      end

        751 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   751");
      end

        752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   752");
      end

        753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   753");
      end

        754 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   754");
      end

        755 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   755");
      end

        756 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   756");
      end

        757 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   757");
      end

        758 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   758");
      end

        759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   759");
      end

        760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   760");
      end

        761 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   761");
      end

        762 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   762");
      end

        763 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   763");
      end

        764 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   764");
      end

        765 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   765");
      end

        766 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   766");
      end

        767 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   767");
      end

        768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   768");
      end

        769 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   769");
      end

        770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   770");
      end

        771 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   771");
      end

        772 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   772");
      end

        773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   773");
      end

        774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   774");
      end

        775 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   775");
      end

        776 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   776");
      end

        777 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   777");
      end

        778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   778");
      end

        779 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   779");
      end

        780 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   780");
      end

        781 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   781");
      end

        782 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   782");
      end

        783 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   783");
      end

        784 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   784");
      end

        785 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   785");
      end

        786 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   786");
      end

        787 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   787");
      end

        788 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   788");
      end

        789 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   789");
      end

        790 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   790");
      end

        791 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   791");
      end

        792 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   792");
      end

        793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   793");
      end

        794 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   794");
      end

        795 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   795");
      end

        796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   796");
      end

        797 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   797");
      end

        798 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   798");
      end

        799 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   799");
      end

        800 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   800");
      end

        801 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   801");
      end

        802 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
         $display("Should not be executed   802");
      end

        803 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   803");
      end

        804 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   804");
      end

        805 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   805");
      end

        806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   806");
      end

        807 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   807");
      end

        808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   808");
      end

        809 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   809");
      end

        810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   810");
      end

        811 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   811");
      end

        812 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   812");
      end

        813 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   813");
      end

        814 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   814");
      end

        815 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   815");
      end

        816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   816");
      end

        817 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   817");
      end

        818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   818");
      end

        819 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   819");
      end

        820 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   820");
      end

        821 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   821");
      end

        822 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   822");
      end

        823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   823");
      end

        824 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   824");
      end

        825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   825");
      end

        826 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   826");
      end

        827 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   827");
      end

        828 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   828");
      end

        829 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   829");
      end

        830 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   830");
      end

        831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   831");
      end

        832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   832");
      end

        833 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   833");
      end

        834 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed   834");
      end

        835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   835");
      end

        836 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed   836");
      end

        837 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   837");
      end

        838 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   838");
      end

        839 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed   839");
      end

        840 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   840");
      end

        841 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   841");
      end

        842 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   842");
      end

        843 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   843");
      end

        844 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   844");
      end

        845 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   845");
      end

        846 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   846");
      end

        847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   847");
      end

        848 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   848");
      end

        849 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   849");
      end

        850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   850");
      end

        851 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   851");
      end

        852 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   852");
      end

        853 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   853");
      end

        854 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   854");
      end

        855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   855");
      end

        856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   856");
      end

        857 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   857");
      end

        858 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   858");
      end

        859 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   859");
      end

        860 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   860");
      end

        861 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   861");
      end

        862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   862");
      end

        863 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   863");
      end

        864 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   864");
      end

        865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   865");
      end

        866 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   866");
      end

        867 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   867");
      end

        868 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   868");
      end

        869 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   869");
      end

        870 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   870");
      end

        871 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   871");
      end

        872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   872");
      end

        873 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   873");
      end

        874 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   874");
      end

        875 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   875");
      end

        876 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   876");
      end

        877 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   877");
      end

        878 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   878");
      end

        879 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   879");
      end

        880 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   880");
      end

        881 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   881");
      end

        882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   882");
      end

        883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   883");
      end

        884 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   884");
      end

        885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   885");
      end

        886 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   886");
      end

        887 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   887");
      end

        888 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   888");
      end

        889 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   889");
      end

        890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   890");
      end

        891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   891");
      end

        892 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   892");
      end

        893 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   893");
      end

        894 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   894");
      end

        895 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   895");
      end

        896 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   896");
      end

        897 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   897");
      end

        898 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   898");
      end

        899 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   899");
      end

        900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   900");
      end

        901 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   901");
      end

        902 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   902");
      end

        903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   903");
      end

        904 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   904");
      end

        905 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   905");
      end

        906 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   906");
      end

        907 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   907");
      end

        908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   908");
      end

        909 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   909");
      end

        910 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   910");
      end

        911 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   911");
      end

        912 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   912");
      end

        913 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   913");
      end

        914 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed   914");
      end

        915 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   915");
      end

        916 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed   916");
      end

        917 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed   917");
      end

        918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   918");
      end

        919 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   919");
      end

        920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   920");
      end

        921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   921");
      end

        922 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   922");
      end

        923 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   923");
      end

        924 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   924");
      end

        925 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed   925");
      end

        926 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   926");
      end

        927 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   927");
      end

        928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   928");
      end

        929 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   929");
      end

        930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   930");
      end

        931 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   931");
      end

        932 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed   932");
      end

        933 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   933");
      end

        934 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   934");
      end

        935 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   935");
      end

        936 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   936");
      end

        937 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   937");
      end

        938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   938");
      end

        939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   939");
      end

        940 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   940");
      end

        941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   941");
      end

        942 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   942");
      end

        943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   943");
      end

        944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   944");
      end

        945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   945");
      end

        946 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   946");
      end

        947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   947");
      end

        948 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   948");
      end

        949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   949");
      end

        950 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   950");
      end

        951 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   951");
      end

        952 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   952");
      end

        953 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   953");
      end

        954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   954");
      end

        955 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   955");
      end

        956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   956");
      end

        957 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   957");
      end

        958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   958");
      end

        959 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed   959");
      end

        960 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed   960");
      end

        961 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   961");
      end

        962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   962");
      end

        963 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed   963");
      end

        964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   964");
      end

        965 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   965");
      end

        966 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   966");
      end

        967 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   967");
      end

        968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   968");
      end

        969 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   969");
      end

        970 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   970");
      end

        971 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   971");
      end

        972 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   972");
      end

        973 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   973");
      end

        974 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   974");
      end

        975 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   975");
      end

        976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   976");
      end

        977 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   977");
      end

        978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   978");
      end

        979 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   979");
      end

        980 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   980");
      end

        981 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   981");
      end

        982 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   982");
      end

        983 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   983");
      end

        984 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed   984");
      end

        985 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   985");
      end

        986 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   986");
      end

        987 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   987");
      end

        988 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   988");
      end

        989 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   989");
      end

        990 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   990");
      end

        991 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed   991");
      end

        992 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   992");
      end

        993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   993");
      end

        994 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   994");
      end

        995 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   995");
      end

        996 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed   996");
      end

        997 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed   997");
      end

        998 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed   998");
      end

        999 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed   999");
      end

       1000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1000");
      end

       1001 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1001");
      end

       1002 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1002");
      end

       1003 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1003");
      end

       1004 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1004");
      end

       1005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1005");
      end

       1006 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1006");
      end

       1007 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1007");
      end

       1008 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1008");
      end

       1009 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1009");
      end

       1010 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1010");
      end

       1011 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1011");
      end

       1012 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1012");
      end

       1013 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1013");
      end

       1014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1014");
      end

       1015 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1015");
      end

       1016 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1016");
      end

       1017 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1017");
      end

       1018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1018");
      end

       1019 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1019");
      end

       1020 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1020");
      end

       1021 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1021");
      end

       1022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1022");
      end

       1023 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1023");
      end

       1024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1024");
      end

       1025 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1025");
      end

       1026 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1026");
      end

       1027 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1027");
      end

       1028 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1028");
      end

       1029 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1029");
      end

       1030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1030");
      end

       1031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1031");
      end

       1032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1032");
      end

       1033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1033");
      end

       1034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1034");
      end

       1035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1035");
      end

       1036 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1036");
      end

       1037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1037");
      end

       1038 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1038");
      end

       1039 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1039");
      end

       1040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1040");
      end

       1041 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1041");
      end

       1042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1042");
      end

       1043 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1043");
      end

       1044 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1044");
      end

       1045 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1045");
      end

       1046 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1046");
      end

       1047 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1047");
      end

       1048 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1048");
      end

       1049 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1049");
      end

       1050 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1050");
      end

       1051 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1051");
      end

       1052 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1052");
      end

       1053 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1053");
      end

       1054 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1054");
      end

       1055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1055");
      end

       1056 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1056");
      end

       1057 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1057");
      end

       1058 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1058");
      end

       1059 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1060;
      end

       1060 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[1]] = 0;
              freedArrays[freedArraysTop] = localMem[1];
              freedArraysTop = freedArraysTop + 1;
              ip = 1061;
      end

       1061 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[476] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[476] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[476]] = 0;
              ip = 1062;
      end

       1062 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1063;
      end

       1063 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[477] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 1064;
      end

       1064 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[477] != 0 ? 1087 : 1065;
      end

       1065 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1065");
      end

       1066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1066");
      end

       1067 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1067");
      end

       1068 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1068");
      end

       1069 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1069");
      end

       1070 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1070");
      end

       1071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1071");
      end

       1072 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1072");
      end

       1073 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1073");
      end

       1074 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1074");
      end

       1075 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1075");
      end

       1076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1076");
      end

       1077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1077");
      end

       1078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1078");
      end

       1079 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1079");
      end

       1080 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1080");
      end

       1081 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1081");
      end

       1082 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1082");
      end

       1083 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1083");
      end

       1084 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1084");
      end

       1085 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1085");
      end

       1086 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1086");
      end

       1087 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1088;
      end

       1088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[485] = heapMem[localMem[477]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 1089;
      end

       1089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[486] = heapMem[localMem[0]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1090;
      end

       1090 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[485] >= localMem[486] ? 1126 : 1091;
      end

       1091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[487] = heapMem[localMem[477]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 1092;
      end

       1092 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[487] != 0 ? 1125 : 1093;
      end

       1093 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[488] = !heapMem[localMem[477]*7 + 6];
              ip = 1094;
      end

       1094 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[488] == 0 ? 1124 : 1095;
      end

       1095 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[489] = heapMem[localMem[477]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1096;
      end

       1096 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[490] = 0; k = arraySizes[localMem[489]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[489] * NArea + i] == 2) localMem[490] = i + 1;
              end
              ip = 1097;
      end

       1097 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[490] == 0 ? 1102 : 1098;
      end

       1098 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1098");
      end

       1099 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1099");
      end

       1100 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1100");
      end

       1101 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1101");
      end

       1102 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 1103;
      end

       1103 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[489]] = localMem[485];
              ip = 1104;
      end

       1104 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[492] = heapMem[localMem[477]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1105;
      end

       1105 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[492]] = localMem[485];
              ip = 1106;
      end

       1106 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[489]];
//$display("AAAAA k=%d  source2=%d", k, 2);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[489] * NArea + i]);
                if (i < k && heapMem[localMem[489] * NArea + i] > 2) j = j + 1;
              end
              localMem[493] = j;
              ip = 1107;
      end

       1107 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[493] != 0 ? 1115 : 1108;
      end

       1108 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[494] = heapMem[localMem[477]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 1109;
      end

       1109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[494]*7 + localMem[485]] = 2;
              updateArrayLength(1, localMem[494], localMem[485]);
              ip = 1110;
      end

       1110 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[495] = heapMem[localMem[477]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 1111;
      end

       1111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[495]*7 + localMem[485]] = 22;
              updateArrayLength(1, localMem[495], localMem[485]);
              ip = 1112;
      end

       1112 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[477]*7 + 0] = localMem[485] + 1;
              updateArrayLength(1, localMem[477], 0);
              ip = 1113;
      end

       1113 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = heapMem[localMem[0]*7 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 1114;
      end

       1114 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 2115;
      end

       1115 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1115");
      end

       1116 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  1116");
      end

       1117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1117");
      end

       1118 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1118");
      end

       1119 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1119");
      end

       1120 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1120");
      end

       1121 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1121");
      end

       1122 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1122");
      end

       1123 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1123");
      end

       1124 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1124");
      end

       1125 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1125");
      end

       1126 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1126");
      end

       1127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1127");
      end

       1128 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1128");
      end

       1129 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1129");
      end

       1130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1130");
      end

       1131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1131");
      end

       1132 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  1132");
      end

       1133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1133");
      end

       1134 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  1134");
      end

       1135 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1135");
      end

       1136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1136");
      end

       1137 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1137");
      end

       1138 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1138");
      end

       1139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1139");
      end

       1140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1140");
      end

       1141 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1141");
      end

       1142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1142");
      end

       1143 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1143");
      end

       1144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1144");
      end

       1145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1145");
      end

       1146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1146");
      end

       1147 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1147");
      end

       1148 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1148");
      end

       1149 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1149");
      end

       1150 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1150");
      end

       1151 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1151");
      end

       1152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1152");
      end

       1153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1153");
      end

       1154 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1154");
      end

       1155 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1155");
      end

       1156 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1156");
      end

       1157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1157");
      end

       1158 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1158");
      end

       1159 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1159");
      end

       1160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1160");
      end

       1161 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1161");
      end

       1162 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1162");
      end

       1163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1163");
      end

       1164 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1164");
      end

       1165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1165");
      end

       1166 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1166");
      end

       1167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1167");
      end

       1168 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1168");
      end

       1169 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1169");
      end

       1170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1170");
      end

       1171 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1171");
      end

       1172 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1172");
      end

       1173 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1173");
      end

       1174 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1174");
      end

       1175 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1175");
      end

       1176 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1176");
      end

       1177 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1177");
      end

       1178 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1178");
      end

       1179 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1179");
      end

       1180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1180");
      end

       1181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1181");
      end

       1182 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1182");
      end

       1183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1183");
      end

       1184 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1184");
      end

       1185 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1185");
      end

       1186 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1186");
      end

       1187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1187");
      end

       1188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1188");
      end

       1189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1189");
      end

       1190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1190");
      end

       1191 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1191");
      end

       1192 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1192");
      end

       1193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1193");
      end

       1194 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1194");
      end

       1195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1195");
      end

       1196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1196");
      end

       1197 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1197");
      end

       1198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1198");
      end

       1199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1199");
      end

       1200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1200");
      end

       1201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1201");
      end

       1202 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1202");
      end

       1203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1203");
      end

       1204 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1204");
      end

       1205 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1205");
      end

       1206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1206");
      end

       1207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1207");
      end

       1208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1208");
      end

       1209 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1209");
      end

       1210 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1210");
      end

       1211 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1211");
      end

       1212 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  1212");
      end

       1213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1213");
      end

       1214 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  1214");
      end

       1215 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1215");
      end

       1216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1216");
      end

       1217 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1217");
      end

       1218 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1218");
      end

       1219 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1219");
      end

       1220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1220");
      end

       1221 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1221");
      end

       1222 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1222");
      end

       1223 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1223");
      end

       1224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1224");
      end

       1225 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1225");
      end

       1226 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1226");
      end

       1227 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1227");
      end

       1228 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1228");
      end

       1229 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1229");
      end

       1230 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1230");
      end

       1231 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1231");
      end

       1232 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1232");
      end

       1233 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1233");
      end

       1234 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1234");
      end

       1235 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1235");
      end

       1236 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1236");
      end

       1237 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1237");
      end

       1238 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1238");
      end

       1239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1239");
      end

       1240 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1240");
      end

       1241 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1241");
      end

       1242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1242");
      end

       1243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1243");
      end

       1244 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1244");
      end

       1245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1245");
      end

       1246 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1246");
      end

       1247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1247");
      end

       1248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1248");
      end

       1249 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1249");
      end

       1250 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1250");
      end

       1251 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1251");
      end

       1252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1252");
      end

       1253 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1253");
      end

       1254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1254");
      end

       1255 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1255");
      end

       1256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1256");
      end

       1257 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1257");
      end

       1258 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1258");
      end

       1259 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1259");
      end

       1260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1260");
      end

       1261 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1261");
      end

       1262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1262");
      end

       1263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1263");
      end

       1264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1264");
      end

       1265 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1265");
      end

       1266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1266");
      end

       1267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1267");
      end

       1268 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1268");
      end

       1269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1269");
      end

       1270 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1270");
      end

       1271 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1271");
      end

       1272 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1272");
      end

       1273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1273");
      end

       1274 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1274");
      end

       1275 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1275");
      end

       1276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1276");
      end

       1277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1277");
      end

       1278 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1278");
      end

       1279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1279");
      end

       1280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1280");
      end

       1281 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1281");
      end

       1282 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1282");
      end

       1283 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1283");
      end

       1284 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1284");
      end

       1285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1285");
      end

       1286 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1286");
      end

       1287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1287");
      end

       1288 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1288");
      end

       1289 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1289");
      end

       1290 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1290");
      end

       1291 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1291");
      end

       1292 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1292");
      end

       1293 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1293");
      end

       1294 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1294");
      end

       1295 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1295");
      end

       1296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1296");
      end

       1297 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1297");
      end

       1298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1298");
      end

       1299 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1299");
      end

       1300 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1300");
      end

       1301 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1301");
      end

       1302 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1302");
      end

       1303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1303");
      end

       1304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1304");
      end

       1305 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1305");
      end

       1306 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1306");
      end

       1307 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1307");
      end

       1308 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1308");
      end

       1309 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1309");
      end

       1310 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1310");
      end

       1311 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1311");
      end

       1312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1312");
      end

       1313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1313");
      end

       1314 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1314");
      end

       1315 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1315");
      end

       1316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1316");
      end

       1317 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1317");
      end

       1318 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1318");
      end

       1319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1319");
      end

       1320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1320");
      end

       1321 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1321");
      end

       1322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1322");
      end

       1323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1323");
      end

       1324 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1324");
      end

       1325 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1325");
      end

       1326 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1326");
      end

       1327 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1327");
      end

       1328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1328");
      end

       1329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1329");
      end

       1330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1330");
      end

       1331 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1331");
      end

       1332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1332");
      end

       1333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1333");
      end

       1334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1334");
      end

       1335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1335");
      end

       1336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1336");
      end

       1337 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1337");
      end

       1338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1338");
      end

       1339 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1339");
      end

       1340 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1340");
      end

       1341 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1341");
      end

       1342 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1342");
      end

       1343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1343");
      end

       1344 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1344");
      end

       1345 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1345");
      end

       1346 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1346");
      end

       1347 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1347");
      end

       1348 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1348");
      end

       1349 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1349");
      end

       1350 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1350");
      end

       1351 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1351");
      end

       1352 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1352");
      end

       1353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1353");
      end

       1354 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1354");
      end

       1355 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1355");
      end

       1356 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1356");
      end

       1357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1357");
      end

       1358 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1358");
      end

       1359 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1359");
      end

       1360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1360");
      end

       1361 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1361");
      end

       1362 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1362");
      end

       1363 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1363");
      end

       1364 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
         $display("Should not be executed  1364");
      end

       1365 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1365");
      end

       1366 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1366");
      end

       1367 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1367");
      end

       1368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1368");
      end

       1369 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1369");
      end

       1370 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1370");
      end

       1371 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1371");
      end

       1372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1372");
      end

       1373 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1373");
      end

       1374 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1374");
      end

       1375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1375");
      end

       1376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1376");
      end

       1377 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1377");
      end

       1378 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  1378");
      end

       1379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1379");
      end

       1380 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  1380");
      end

       1381 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1381");
      end

       1382 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1382");
      end

       1383 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1383");
      end

       1384 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1384");
      end

       1385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1385");
      end

       1386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1386");
      end

       1387 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1387");
      end

       1388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1388");
      end

       1389 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1389");
      end

       1390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1390");
      end

       1391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1391");
      end

       1392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1392");
      end

       1393 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1393");
      end

       1394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1394");
      end

       1395 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1395");
      end

       1396 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1396");
      end

       1397 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1397");
      end

       1398 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1398");
      end

       1399 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1399");
      end

       1400 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1400");
      end

       1401 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1401");
      end

       1402 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1402");
      end

       1403 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1403");
      end

       1404 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1404");
      end

       1405 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1405");
      end

       1406 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1406");
      end

       1407 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1407");
      end

       1408 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1408");
      end

       1409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1409");
      end

       1410 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1410");
      end

       1411 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1411");
      end

       1412 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1412");
      end

       1413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1413");
      end

       1414 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1414");
      end

       1415 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1415");
      end

       1416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1416");
      end

       1417 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1417");
      end

       1418 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1418");
      end

       1419 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1419");
      end

       1420 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1420");
      end

       1421 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1421");
      end

       1422 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1422");
      end

       1423 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1423");
      end

       1424 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1424");
      end

       1425 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1425");
      end

       1426 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1426");
      end

       1427 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1427");
      end

       1428 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1428");
      end

       1429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1429");
      end

       1430 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1430");
      end

       1431 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1431");
      end

       1432 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1432");
      end

       1433 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1433");
      end

       1434 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1434");
      end

       1435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1435");
      end

       1436 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1436");
      end

       1437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1437");
      end

       1438 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1438");
      end

       1439 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1439");
      end

       1440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1440");
      end

       1441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1441");
      end

       1442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1442");
      end

       1443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1443");
      end

       1444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1444");
      end

       1445 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1445");
      end

       1446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1446");
      end

       1447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1447");
      end

       1448 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1448");
      end

       1449 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1449");
      end

       1450 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1450");
      end

       1451 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1451");
      end

       1452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1452");
      end

       1453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1453");
      end

       1454 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1454");
      end

       1455 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1455");
      end

       1456 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1456");
      end

       1457 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1457");
      end

       1458 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  1458");
      end

       1459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1459");
      end

       1460 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  1460");
      end

       1461 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1461");
      end

       1462 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1462");
      end

       1463 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1463");
      end

       1464 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1464");
      end

       1465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1465");
      end

       1466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1466");
      end

       1467 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1467");
      end

       1468 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1468");
      end

       1469 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1469");
      end

       1470 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1470");
      end

       1471 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1471");
      end

       1472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1472");
      end

       1473 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1473");
      end

       1474 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1474");
      end

       1475 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1475");
      end

       1476 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1476");
      end

       1477 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1477");
      end

       1478 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1478");
      end

       1479 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1479");
      end

       1480 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1480");
      end

       1481 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1481");
      end

       1482 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1482");
      end

       1483 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1483");
      end

       1484 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1484");
      end

       1485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1485");
      end

       1486 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1486");
      end

       1487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1487");
      end

       1488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1488");
      end

       1489 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1489");
      end

       1490 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1490");
      end

       1491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1491");
      end

       1492 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1492");
      end

       1493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1493");
      end

       1494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1494");
      end

       1495 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1495");
      end

       1496 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1496");
      end

       1497 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1497");
      end

       1498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1498");
      end

       1499 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1499");
      end

       1500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1500");
      end

       1501 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1501");
      end

       1502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1502");
      end

       1503 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1503");
      end

       1504 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1504");
      end

       1505 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1505");
      end

       1506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1506");
      end

       1507 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1507");
      end

       1508 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1508");
      end

       1509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1509");
      end

       1510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1510");
      end

       1511 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1511");
      end

       1512 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1512");
      end

       1513 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1513");
      end

       1514 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1514");
      end

       1515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1515");
      end

       1516 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1516");
      end

       1517 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1517");
      end

       1518 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1518");
      end

       1519 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1519");
      end

       1520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1520");
      end

       1521 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1521");
      end

       1522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1522");
      end

       1523 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1523");
      end

       1524 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1524");
      end

       1525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1525");
      end

       1526 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1526");
      end

       1527 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1527");
      end

       1528 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1528");
      end

       1529 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1529");
      end

       1530 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1530");
      end

       1531 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1531");
      end

       1532 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1532");
      end

       1533 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1533");
      end

       1534 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1534");
      end

       1535 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1535");
      end

       1536 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1536");
      end

       1537 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1537");
      end

       1538 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1538");
      end

       1539 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1539");
      end

       1540 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1540");
      end

       1541 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1541");
      end

       1542 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1542");
      end

       1543 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1543");
      end

       1544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1544");
      end

       1545 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1545");
      end

       1546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1546");
      end

       1547 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1547");
      end

       1548 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1548");
      end

       1549 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1549");
      end

       1550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1550");
      end

       1551 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1551");
      end

       1552 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1552");
      end

       1553 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1553");
      end

       1554 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1554");
      end

       1555 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1555");
      end

       1556 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1556");
      end

       1557 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1557");
      end

       1558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1558");
      end

       1559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1559");
      end

       1560 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1560");
      end

       1561 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1561");
      end

       1562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1562");
      end

       1563 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1563");
      end

       1564 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1564");
      end

       1565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1565");
      end

       1566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1566");
      end

       1567 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1567");
      end

       1568 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1568");
      end

       1569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1569");
      end

       1570 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1570");
      end

       1571 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1571");
      end

       1572 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1572");
      end

       1573 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1573");
      end

       1574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1574");
      end

       1575 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1575");
      end

       1576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1576");
      end

       1577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1577");
      end

       1578 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1578");
      end

       1579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1579");
      end

       1580 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1580");
      end

       1581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1581");
      end

       1582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1582");
      end

       1583 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1583");
      end

       1584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1584");
      end

       1585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1585");
      end

       1586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1586");
      end

       1587 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1587");
      end

       1588 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1588");
      end

       1589 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1589");
      end

       1590 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1590");
      end

       1591 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1591");
      end

       1592 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1592");
      end

       1593 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1593");
      end

       1594 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1594");
      end

       1595 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1595");
      end

       1596 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1596");
      end

       1597 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1597");
      end

       1598 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1598");
      end

       1599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1599");
      end

       1600 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1600");
      end

       1601 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1601");
      end

       1602 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1602");
      end

       1603 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1603");
      end

       1604 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1604");
      end

       1605 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1605");
      end

       1606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1606");
      end

       1607 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  1607");
      end

       1608 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1608");
      end

       1609 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1609");
      end

       1610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1610");
      end

       1611 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1611");
      end

       1612 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1612");
      end

       1613 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1613");
      end

       1614 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  1614");
      end

       1615 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1615");
      end

       1616 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1616");
      end

       1617 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1617");
      end

       1618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1618");
      end

       1619 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1619");
      end

       1620 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1620");
      end

       1621 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1621");
      end

       1622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1622");
      end

       1623 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1623");
      end

       1624 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1624");
      end

       1625 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1625");
      end

       1626 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1626");
      end

       1627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1627");
      end

       1628 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  1628");
      end

       1629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1629");
      end

       1630 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  1630");
      end

       1631 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1631");
      end

       1632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1632");
      end

       1633 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1633");
      end

       1634 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1634");
      end

       1635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1635");
      end

       1636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1636");
      end

       1637 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1637");
      end

       1638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1638");
      end

       1639 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1639");
      end

       1640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1640");
      end

       1641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1641");
      end

       1642 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1642");
      end

       1643 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1643");
      end

       1644 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1644");
      end

       1645 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1645");
      end

       1646 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1646");
      end

       1647 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1647");
      end

       1648 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1648");
      end

       1649 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1649");
      end

       1650 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1650");
      end

       1651 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1651");
      end

       1652 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1652");
      end

       1653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1653");
      end

       1654 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1654");
      end

       1655 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1655");
      end

       1656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1656");
      end

       1657 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1657");
      end

       1658 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1658");
      end

       1659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1659");
      end

       1660 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1660");
      end

       1661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1661");
      end

       1662 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1662");
      end

       1663 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1663");
      end

       1664 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1664");
      end

       1665 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1665");
      end

       1666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1666");
      end

       1667 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1667");
      end

       1668 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1668");
      end

       1669 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1669");
      end

       1670 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1670");
      end

       1671 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1671");
      end

       1672 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1672");
      end

       1673 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1673");
      end

       1674 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1674");
      end

       1675 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1675");
      end

       1676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1676");
      end

       1677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1677");
      end

       1678 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1678");
      end

       1679 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1679");
      end

       1680 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1680");
      end

       1681 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1681");
      end

       1682 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1682");
      end

       1683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1683");
      end

       1684 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1684");
      end

       1685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1685");
      end

       1686 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1686");
      end

       1687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1687");
      end

       1688 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1688");
      end

       1689 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1689");
      end

       1690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1690");
      end

       1691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1691");
      end

       1692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1692");
      end

       1693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1693");
      end

       1694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1694");
      end

       1695 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1695");
      end

       1696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1696");
      end

       1697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1697");
      end

       1698 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1698");
      end

       1699 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1699");
      end

       1700 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1700");
      end

       1701 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1701");
      end

       1702 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1702");
      end

       1703 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1703");
      end

       1704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1704");
      end

       1705 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1705");
      end

       1706 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1706");
      end

       1707 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1707");
      end

       1708 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  1708");
      end

       1709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1709");
      end

       1710 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  1710");
      end

       1711 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1711");
      end

       1712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1712");
      end

       1713 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1713");
      end

       1714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1714");
      end

       1715 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1715");
      end

       1716 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1716");
      end

       1717 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1717");
      end

       1718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1718");
      end

       1719 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1719");
      end

       1720 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1720");
      end

       1721 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1721");
      end

       1722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1722");
      end

       1723 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1723");
      end

       1724 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1724");
      end

       1725 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1725");
      end

       1726 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1726");
      end

       1727 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1727");
      end

       1728 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1728");
      end

       1729 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1729");
      end

       1730 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1730");
      end

       1731 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1731");
      end

       1732 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1732");
      end

       1733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1733");
      end

       1734 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1734");
      end

       1735 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1735");
      end

       1736 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1736");
      end

       1737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1737");
      end

       1738 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1738");
      end

       1739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1739");
      end

       1740 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1740");
      end

       1741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1741");
      end

       1742 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1742");
      end

       1743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1743");
      end

       1744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1744");
      end

       1745 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1745");
      end

       1746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1746");
      end

       1747 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1747");
      end

       1748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1748");
      end

       1749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1749");
      end

       1750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1750");
      end

       1751 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1751");
      end

       1752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1752");
      end

       1753 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1753");
      end

       1754 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1754");
      end

       1755 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1755");
      end

       1756 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1756");
      end

       1757 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1757");
      end

       1758 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1758");
      end

       1759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1759");
      end

       1760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1760");
      end

       1761 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1761");
      end

       1762 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1762");
      end

       1763 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1763");
      end

       1764 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1764");
      end

       1765 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1765");
      end

       1766 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1766");
      end

       1767 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1767");
      end

       1768 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1768");
      end

       1769 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1769");
      end

       1770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1770");
      end

       1771 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1771");
      end

       1772 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1772");
      end

       1773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1773");
      end

       1774 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1774");
      end

       1775 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1775");
      end

       1776 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1776");
      end

       1777 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1777");
      end

       1778 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1778");
      end

       1779 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1779");
      end

       1780 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1780");
      end

       1781 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1781");
      end

       1782 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1782");
      end

       1783 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1783");
      end

       1784 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1784");
      end

       1785 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1785");
      end

       1786 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1786");
      end

       1787 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1787");
      end

       1788 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1788");
      end

       1789 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1789");
      end

       1790 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1790");
      end

       1791 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1791");
      end

       1792 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1792");
      end

       1793 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1793");
      end

       1794 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1794");
      end

       1795 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1795");
      end

       1796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1796");
      end

       1797 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1797");
      end

       1798 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1798");
      end

       1799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1799");
      end

       1800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1800");
      end

       1801 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1801");
      end

       1802 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1802");
      end

       1803 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1803");
      end

       1804 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1804");
      end

       1805 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1805");
      end

       1806 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1806");
      end

       1807 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1807");
      end

       1808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1808");
      end

       1809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1809");
      end

       1810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1810");
      end

       1811 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1811");
      end

       1812 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1812");
      end

       1813 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1813");
      end

       1814 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1814");
      end

       1815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1815");
      end

       1816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1816");
      end

       1817 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1817");
      end

       1818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1818");
      end

       1819 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1819");
      end

       1820 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1820");
      end

       1821 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1821");
      end

       1822 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1822");
      end

       1823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1823");
      end

       1824 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1824");
      end

       1825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1825");
      end

       1826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1826");
      end

       1827 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1827");
      end

       1828 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1828");
      end

       1829 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1829");
      end

       1830 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1830");
      end

       1831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1831");
      end

       1832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1832");
      end

       1833 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1833");
      end

       1834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1834");
      end

       1835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1835");
      end

       1836 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1836");
      end

       1837 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1837");
      end

       1838 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1838");
      end

       1839 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1839");
      end

       1840 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1840");
      end

       1841 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1841");
      end

       1842 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1842");
      end

       1843 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1843");
      end

       1844 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1844");
      end

       1845 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1845");
      end

       1846 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1846");
      end

       1847 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1847");
      end

       1848 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1848");
      end

       1849 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1849");
      end

       1850 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1850");
      end

       1851 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1851");
      end

       1852 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1852");
      end

       1853 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1853");
      end

       1854 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1854");
      end

       1855 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1855");
      end

       1856 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1856");
      end

       1857 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1857");
      end

       1858 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
         $display("Should not be executed  1858");
      end

       1859 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1859");
      end

       1860 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1860");
      end

       1861 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1861");
      end

       1862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1862");
      end

       1863 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1863");
      end

       1864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1864");
      end

       1865 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1865");
      end

       1866 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1866");
      end

       1867 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1867");
      end

       1868 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1868");
      end

       1869 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1869");
      end

       1870 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1870");
      end

       1871 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1871");
      end

       1872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1872");
      end

       1873 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1873");
      end

       1874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1874");
      end

       1875 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1875");
      end

       1876 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1876");
      end

       1877 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1877");
      end

       1878 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1878");
      end

       1879 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1879");
      end

       1880 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1880");
      end

       1881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1881");
      end

       1882 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1882");
      end

       1883 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1883");
      end

       1884 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1884");
      end

       1885 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1885");
      end

       1886 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1886");
      end

       1887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1887");
      end

       1888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1888");
      end

       1889 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1889");
      end

       1890 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  1890");
      end

       1891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1891");
      end

       1892 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  1892");
      end

       1893 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1893");
      end

       1894 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1894");
      end

       1895 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  1895");
      end

       1896 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1896");
      end

       1897 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1897");
      end

       1898 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1898");
      end

       1899 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1899");
      end

       1900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1900");
      end

       1901 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1901");
      end

       1902 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1902");
      end

       1903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1903");
      end

       1904 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1904");
      end

       1905 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1905");
      end

       1906 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1906");
      end

       1907 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  1907");
      end

       1908 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1908");
      end

       1909 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1909");
      end

       1910 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1910");
      end

       1911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1911");
      end

       1912 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1912");
      end

       1913 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1913");
      end

       1914 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1914");
      end

       1915 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1915");
      end

       1916 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1916");
      end

       1917 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1917");
      end

       1918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1918");
      end

       1919 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1919");
      end

       1920 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1920");
      end

       1921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1921");
      end

       1922 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1922");
      end

       1923 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1923");
      end

       1924 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1924");
      end

       1925 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1925");
      end

       1926 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1926");
      end

       1927 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  1927");
      end

       1928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1928");
      end

       1929 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1929");
      end

       1930 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1930");
      end

       1931 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1931");
      end

       1932 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1932");
      end

       1933 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1933");
      end

       1934 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1934");
      end

       1935 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1935");
      end

       1936 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1936");
      end

       1937 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1937");
      end

       1938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1938");
      end

       1939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1939");
      end

       1940 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1940");
      end

       1941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1941");
      end

       1942 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1942");
      end

       1943 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  1943");
      end

       1944 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1944");
      end

       1945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1945");
      end

       1946 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1946");
      end

       1947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1947");
      end

       1948 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1948");
      end

       1949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1949");
      end

       1950 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  1950");
      end

       1951 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1951");
      end

       1952 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1952");
      end

       1953 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1953");
      end

       1954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1954");
      end

       1955 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1955");
      end

       1956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1956");
      end

       1957 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1957");
      end

       1958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1958");
      end

       1959 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1959");
      end

       1960 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1960");
      end

       1961 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1961");
      end

       1962 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1962");
      end

       1963 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1963");
      end

       1964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1964");
      end

       1965 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1965");
      end

       1966 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1966");
      end

       1967 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1967");
      end

       1968 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1968");
      end

       1969 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1969");
      end

       1970 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  1970");
      end

       1971 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1971");
      end

       1972 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  1972");
      end

       1973 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  1973");
      end

       1974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1974");
      end

       1975 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1975");
      end

       1976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1976");
      end

       1977 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1977");
      end

       1978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1978");
      end

       1979 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1979");
      end

       1980 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1980");
      end

       1981 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  1981");
      end

       1982 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1982");
      end

       1983 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1983");
      end

       1984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1984");
      end

       1985 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1985");
      end

       1986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1986");
      end

       1987 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1987");
      end

       1988 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  1988");
      end

       1989 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  1989");
      end

       1990 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  1990");
      end

       1991 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1991");
      end

       1992 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  1992");
      end

       1993 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1993");
      end

       1994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1994");
      end

       1995 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1995");
      end

       1996 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1996");
      end

       1997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1997");
      end

       1998 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  1998");
      end

       1999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  1999");
      end

       2000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2000");
      end

       2001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2001");
      end

       2002 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2002");
      end

       2003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2003");
      end

       2004 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2004");
      end

       2005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2005");
      end

       2006 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2006");
      end

       2007 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2007");
      end

       2008 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2008");
      end

       2009 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2009");
      end

       2010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2010");
      end

       2011 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2011");
      end

       2012 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2012");
      end

       2013 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2013");
      end

       2014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2014");
      end

       2015 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2015");
      end

       2016 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2016");
      end

       2017 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2017");
      end

       2018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2018");
      end

       2019 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2019");
      end

       2020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2020");
      end

       2021 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2021");
      end

       2022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2022");
      end

       2023 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2023");
      end

       2024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2024");
      end

       2025 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2025");
      end

       2026 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2026");
      end

       2027 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2027");
      end

       2028 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2028");
      end

       2029 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2029");
      end

       2030 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2030");
      end

       2031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2031");
      end

       2032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2032");
      end

       2033 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2033");
      end

       2034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2034");
      end

       2035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2035");
      end

       2036 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2036");
      end

       2037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2037");
      end

       2038 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2038");
      end

       2039 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2039");
      end

       2040 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2040");
      end

       2041 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2041");
      end

       2042 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2042");
      end

       2043 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2043");
      end

       2044 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2044");
      end

       2045 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2045");
      end

       2046 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2046");
      end

       2047 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2047");
      end

       2048 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2048");
      end

       2049 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2049");
      end

       2050 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2050");
      end

       2051 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2051");
      end

       2052 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2052");
      end

       2053 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2053");
      end

       2054 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2054");
      end

       2055 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2055");
      end

       2056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2056");
      end

       2057 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2057");
      end

       2058 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2058");
      end

       2059 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2059");
      end

       2060 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2060");
      end

       2061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2061");
      end

       2062 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2062");
      end

       2063 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2063");
      end

       2064 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2064");
      end

       2065 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2065");
      end

       2066 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2066");
      end

       2067 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2067");
      end

       2068 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2068");
      end

       2069 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2069");
      end

       2070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2070");
      end

       2071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2071");
      end

       2072 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2072");
      end

       2073 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2073");
      end

       2074 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2074");
      end

       2075 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2075");
      end

       2076 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2076");
      end

       2077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2077");
      end

       2078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2078");
      end

       2079 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2079");
      end

       2080 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2080");
      end

       2081 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2081");
      end

       2082 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2082");
      end

       2083 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2083");
      end

       2084 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2084");
      end

       2085 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2085");
      end

       2086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2086");
      end

       2087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2087");
      end

       2088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2088");
      end

       2089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2089");
      end

       2090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2090");
      end

       2091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2091");
      end

       2092 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2092");
      end

       2093 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2093");
      end

       2094 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2094");
      end

       2095 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2095");
      end

       2096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2096");
      end

       2097 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2097");
      end

       2098 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2098");
      end

       2099 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2099");
      end

       2100 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2100");
      end

       2101 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2101");
      end

       2102 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2102");
      end

       2103 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2103");
      end

       2104 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2104");
      end

       2105 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2105");
      end

       2106 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2106");
      end

       2107 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2107");
      end

       2108 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2108");
      end

       2109 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2109");
      end

       2110 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2110");
      end

       2111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2111");
      end

       2112 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2112");
      end

       2113 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2113");
      end

       2114 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2114");
      end

       2115 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2116;
      end

       2116 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[476]] = 0;
              freedArrays[freedArraysTop] = localMem[476];
              freedArraysTop = freedArraysTop + 1;
              ip = 2117;
      end

       2117 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[951] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[951] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[951]] = 0;
              ip = 2118;
      end

       2118 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2119;
      end

       2119 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[952] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 2120;
      end

       2120 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[952] != 0 ? 2143 : 2121;
      end

       2121 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2121");
      end

       2122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2122");
      end

       2123 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2123");
      end

       2124 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2124");
      end

       2125 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2125");
      end

       2126 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2126");
      end

       2127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2127");
      end

       2128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2128");
      end

       2129 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2129");
      end

       2130 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2130");
      end

       2131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2131");
      end

       2132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2132");
      end

       2133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2133");
      end

       2134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2134");
      end

       2135 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2135");
      end

       2136 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2136");
      end

       2137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2137");
      end

       2138 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2138");
      end

       2139 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2139");
      end

       2140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2140");
      end

       2141 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2141");
      end

       2142 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2142");
      end

       2143 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2144;
      end

       2144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[960] = heapMem[localMem[952]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 2145;
      end

       2145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[961] = heapMem[localMem[0]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2146;
      end

       2146 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[960] >= localMem[961] ? 2182 : 2147;
      end

       2147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[962] = heapMem[localMem[952]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 2148;
      end

       2148 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[962] != 0 ? 2181 : 2149;
      end

       2149 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[963] = !heapMem[localMem[952]*7 + 6];
              ip = 2150;
      end

       2150 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[963] == 0 ? 2180 : 2151;
      end

       2151 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[964] = heapMem[localMem[952]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2152;
      end

       2152 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
              localMem[965] = 0; k = arraySizes[localMem[964]];
              for(i = 0; i < NArea; i = i + 1) begin
                if (i < k && heapMem[localMem[964] * NArea + i] == 3) localMem[965] = i + 1;
              end
              ip = 2153;
      end

       2153 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[965] == 0 ? 2158 : 2154;
      end

       2154 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2154");
      end

       2155 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2155");
      end

       2156 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2156");
      end

       2157 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2157");
      end

       2158 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 2159;
      end

       2159 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[964]] = localMem[960];
              ip = 2160;
      end

       2160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[967] = heapMem[localMem[952]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2161;
      end

       2161 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[967]] = localMem[960];
              ip = 2162;
      end

       2162 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
              j = 0; k = arraySizes[localMem[964]];
//$display("AAAAA k=%d  source2=%d", k, 3);
              for(i = 0; i < NArea; i = i + 1) begin
//$display("AAAAA i=%d  value=%d", i, heapMem[localMem[964] * NArea + i]);
                if (i < k && heapMem[localMem[964] * NArea + i] > 3) j = j + 1;
              end
              localMem[968] = j;
              ip = 2163;
      end

       2163 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[968] != 0 ? 2171 : 2164;
      end

       2164 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[969] = heapMem[localMem[952]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 2165;
      end

       2165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[969]*7 + localMem[960]] = 3;
              updateArrayLength(1, localMem[969], localMem[960]);
              ip = 2166;
      end

       2166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[970] = heapMem[localMem[952]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 2167;
      end

       2167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[970]*7 + localMem[960]] = 33;
              updateArrayLength(1, localMem[970], localMem[960]);
              ip = 2168;
      end

       2168 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[952]*7 + 0] = localMem[960] + 1;
              updateArrayLength(1, localMem[952], 0);
              ip = 2169;
      end

       2169 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = heapMem[localMem[0]*7 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 2170;
      end

       2170 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3171;
      end

       2171 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2171");
      end

       2172 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  2172");
      end

       2173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2173");
      end

       2174 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2174");
      end

       2175 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2175");
      end

       2176 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2176");
      end

       2177 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2177");
      end

       2178 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2178");
      end

       2179 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2179");
      end

       2180 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2180");
      end

       2181 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2181");
      end

       2182 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2182");
      end

       2183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2183");
      end

       2184 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2184");
      end

       2185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2185");
      end

       2186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2186");
      end

       2187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2187");
      end

       2188 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  2188");
      end

       2189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2189");
      end

       2190 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  2190");
      end

       2191 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2191");
      end

       2192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2192");
      end

       2193 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2193");
      end

       2194 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2194");
      end

       2195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2195");
      end

       2196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2196");
      end

       2197 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2197");
      end

       2198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2198");
      end

       2199 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2199");
      end

       2200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2200");
      end

       2201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2201");
      end

       2202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2202");
      end

       2203 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2203");
      end

       2204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2204");
      end

       2205 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2205");
      end

       2206 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2206");
      end

       2207 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2207");
      end

       2208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2208");
      end

       2209 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2209");
      end

       2210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2210");
      end

       2211 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2211");
      end

       2212 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2212");
      end

       2213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2213");
      end

       2214 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2214");
      end

       2215 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2215");
      end

       2216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2216");
      end

       2217 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2217");
      end

       2218 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2218");
      end

       2219 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2219");
      end

       2220 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2220");
      end

       2221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2221");
      end

       2222 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2222");
      end

       2223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2223");
      end

       2224 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2224");
      end

       2225 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2225");
      end

       2226 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2226");
      end

       2227 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2227");
      end

       2228 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2228");
      end

       2229 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2229");
      end

       2230 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2230");
      end

       2231 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2231");
      end

       2232 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2232");
      end

       2233 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2233");
      end

       2234 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2234");
      end

       2235 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2235");
      end

       2236 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2236");
      end

       2237 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2237");
      end

       2238 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2238");
      end

       2239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2239");
      end

       2240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2240");
      end

       2241 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2241");
      end

       2242 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2242");
      end

       2243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2243");
      end

       2244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2244");
      end

       2245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2245");
      end

       2246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2246");
      end

       2247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2247");
      end

       2248 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2248");
      end

       2249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2249");
      end

       2250 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2250");
      end

       2251 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2251");
      end

       2252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2252");
      end

       2253 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2253");
      end

       2254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2254");
      end

       2255 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2255");
      end

       2256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2256");
      end

       2257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2257");
      end

       2258 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2258");
      end

       2259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2259");
      end

       2260 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2260");
      end

       2261 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2261");
      end

       2262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2262");
      end

       2263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2263");
      end

       2264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2264");
      end

       2265 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2265");
      end

       2266 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2266");
      end

       2267 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2267");
      end

       2268 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  2268");
      end

       2269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2269");
      end

       2270 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  2270");
      end

       2271 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2271");
      end

       2272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2272");
      end

       2273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2273");
      end

       2274 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2274");
      end

       2275 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2275");
      end

       2276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2276");
      end

       2277 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2277");
      end

       2278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2278");
      end

       2279 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2279");
      end

       2280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2280");
      end

       2281 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2281");
      end

       2282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2282");
      end

       2283 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2283");
      end

       2284 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2284");
      end

       2285 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2285");
      end

       2286 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2286");
      end

       2287 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2287");
      end

       2288 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2288");
      end

       2289 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2289");
      end

       2290 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2290");
      end

       2291 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2291");
      end

       2292 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2292");
      end

       2293 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2293");
      end

       2294 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2294");
      end

       2295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2295");
      end

       2296 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2296");
      end

       2297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2297");
      end

       2298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2298");
      end

       2299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2299");
      end

       2300 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2300");
      end

       2301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2301");
      end

       2302 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2302");
      end

       2303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2303");
      end

       2304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2304");
      end

       2305 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2305");
      end

       2306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2306");
      end

       2307 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2307");
      end

       2308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2308");
      end

       2309 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2309");
      end

       2310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2310");
      end

       2311 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2311");
      end

       2312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2312");
      end

       2313 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2313");
      end

       2314 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2314");
      end

       2315 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2315");
      end

       2316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2316");
      end

       2317 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2317");
      end

       2318 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2318");
      end

       2319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2319");
      end

       2320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2320");
      end

       2321 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2321");
      end

       2322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2322");
      end

       2323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2323");
      end

       2324 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2324");
      end

       2325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2325");
      end

       2326 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2326");
      end

       2327 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2327");
      end

       2328 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2328");
      end

       2329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2329");
      end

       2330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2330");
      end

       2331 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2331");
      end

       2332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2332");
      end

       2333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2333");
      end

       2334 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2334");
      end

       2335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2335");
      end

       2336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2336");
      end

       2337 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2337");
      end

       2338 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2338");
      end

       2339 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2339");
      end

       2340 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2340");
      end

       2341 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2341");
      end

       2342 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2342");
      end

       2343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2343");
      end

       2344 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2344");
      end

       2345 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2345");
      end

       2346 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2346");
      end

       2347 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2347");
      end

       2348 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2348");
      end

       2349 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2349");
      end

       2350 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2350");
      end

       2351 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2351");
      end

       2352 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2352");
      end

       2353 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2353");
      end

       2354 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2354");
      end

       2355 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2355");
      end

       2356 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2356");
      end

       2357 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2357");
      end

       2358 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2358");
      end

       2359 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2359");
      end

       2360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2360");
      end

       2361 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2361");
      end

       2362 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2362");
      end

       2363 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2363");
      end

       2364 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2364");
      end

       2365 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2365");
      end

       2366 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2366");
      end

       2367 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2367");
      end

       2368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2368");
      end

       2369 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2369");
      end

       2370 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2370");
      end

       2371 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2371");
      end

       2372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2372");
      end

       2373 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2373");
      end

       2374 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2374");
      end

       2375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2375");
      end

       2376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2376");
      end

       2377 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2377");
      end

       2378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2378");
      end

       2379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2379");
      end

       2380 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2380");
      end

       2381 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2381");
      end

       2382 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2382");
      end

       2383 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2383");
      end

       2384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2384");
      end

       2385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2385");
      end

       2386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2386");
      end

       2387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2387");
      end

       2388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2388");
      end

       2389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2389");
      end

       2390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2390");
      end

       2391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2391");
      end

       2392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2392");
      end

       2393 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2393");
      end

       2394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2394");
      end

       2395 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2395");
      end

       2396 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2396");
      end

       2397 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2397");
      end

       2398 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2398");
      end

       2399 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2399");
      end

       2400 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2400");
      end

       2401 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2401");
      end

       2402 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2402");
      end

       2403 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2403");
      end

       2404 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2404");
      end

       2405 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2405");
      end

       2406 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2406");
      end

       2407 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2407");
      end

       2408 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2408");
      end

       2409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2409");
      end

       2410 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2410");
      end

       2411 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2411");
      end

       2412 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2412");
      end

       2413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2413");
      end

       2414 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2414");
      end

       2415 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2415");
      end

       2416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2416");
      end

       2417 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2417");
      end

       2418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2418");
      end

       2419 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2419");
      end

       2420 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
         $display("Should not be executed  2420");
      end

       2421 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2421");
      end

       2422 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2422");
      end

       2423 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2423");
      end

       2424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2424");
      end

       2425 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2425");
      end

       2426 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2426");
      end

       2427 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2427");
      end

       2428 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2428");
      end

       2429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2429");
      end

       2430 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2430");
      end

       2431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2431");
      end

       2432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2432");
      end

       2433 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2433");
      end

       2434 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  2434");
      end

       2435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2435");
      end

       2436 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  2436");
      end

       2437 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2437");
      end

       2438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2438");
      end

       2439 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2439");
      end

       2440 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2440");
      end

       2441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2441");
      end

       2442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2442");
      end

       2443 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2443");
      end

       2444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2444");
      end

       2445 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2445");
      end

       2446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2446");
      end

       2447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2447");
      end

       2448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2448");
      end

       2449 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2449");
      end

       2450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2450");
      end

       2451 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2451");
      end

       2452 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2452");
      end

       2453 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2453");
      end

       2454 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2454");
      end

       2455 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2455");
      end

       2456 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2456");
      end

       2457 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2457");
      end

       2458 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2458");
      end

       2459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2459");
      end

       2460 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2460");
      end

       2461 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2461");
      end

       2462 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2462");
      end

       2463 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2463");
      end

       2464 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2464");
      end

       2465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2465");
      end

       2466 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2466");
      end

       2467 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2467");
      end

       2468 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2468");
      end

       2469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2469");
      end

       2470 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2470");
      end

       2471 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2471");
      end

       2472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2472");
      end

       2473 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2473");
      end

       2474 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2474");
      end

       2475 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2475");
      end

       2476 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2476");
      end

       2477 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2477");
      end

       2478 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2478");
      end

       2479 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2479");
      end

       2480 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2480");
      end

       2481 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2481");
      end

       2482 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2482");
      end

       2483 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2483");
      end

       2484 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2484");
      end

       2485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2485");
      end

       2486 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2486");
      end

       2487 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2487");
      end

       2488 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2488");
      end

       2489 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2489");
      end

       2490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2490");
      end

       2491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2491");
      end

       2492 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2492");
      end

       2493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2493");
      end

       2494 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2494");
      end

       2495 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2495");
      end

       2496 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2496");
      end

       2497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2497");
      end

       2498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2498");
      end

       2499 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2499");
      end

       2500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2500");
      end

       2501 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2501");
      end

       2502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2502");
      end

       2503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2503");
      end

       2504 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2504");
      end

       2505 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2505");
      end

       2506 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2506");
      end

       2507 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2507");
      end

       2508 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2508");
      end

       2509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2509");
      end

       2510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2510");
      end

       2511 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2511");
      end

       2512 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2512");
      end

       2513 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2513");
      end

       2514 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  2514");
      end

       2515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2515");
      end

       2516 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  2516");
      end

       2517 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2517");
      end

       2518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2518");
      end

       2519 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2519");
      end

       2520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2520");
      end

       2521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2521");
      end

       2522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2522");
      end

       2523 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2523");
      end

       2524 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2524");
      end

       2525 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2525");
      end

       2526 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2526");
      end

       2527 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2527");
      end

       2528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2528");
      end

       2529 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2529");
      end

       2530 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2530");
      end

       2531 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2531");
      end

       2532 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2532");
      end

       2533 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2533");
      end

       2534 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2534");
      end

       2535 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2535");
      end

       2536 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2536");
      end

       2537 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2537");
      end

       2538 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2538");
      end

       2539 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2539");
      end

       2540 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2540");
      end

       2541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2541");
      end

       2542 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2542");
      end

       2543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2543");
      end

       2544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2544");
      end

       2545 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2545");
      end

       2546 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2546");
      end

       2547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2547");
      end

       2548 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2548");
      end

       2549 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2549");
      end

       2550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2550");
      end

       2551 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2551");
      end

       2552 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2552");
      end

       2553 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2553");
      end

       2554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2554");
      end

       2555 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2555");
      end

       2556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2556");
      end

       2557 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2557");
      end

       2558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2558");
      end

       2559 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2559");
      end

       2560 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2560");
      end

       2561 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2561");
      end

       2562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2562");
      end

       2563 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2563");
      end

       2564 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2564");
      end

       2565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2565");
      end

       2566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2566");
      end

       2567 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2567");
      end

       2568 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2568");
      end

       2569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2569");
      end

       2570 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2570");
      end

       2571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2571");
      end

       2572 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2572");
      end

       2573 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2573");
      end

       2574 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2574");
      end

       2575 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2575");
      end

       2576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2576");
      end

       2577 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2577");
      end

       2578 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2578");
      end

       2579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2579");
      end

       2580 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2580");
      end

       2581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2581");
      end

       2582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2582");
      end

       2583 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2583");
      end

       2584 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2584");
      end

       2585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2585");
      end

       2586 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2586");
      end

       2587 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2587");
      end

       2588 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2588");
      end

       2589 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2589");
      end

       2590 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2590");
      end

       2591 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2591");
      end

       2592 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2592");
      end

       2593 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2593");
      end

       2594 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2594");
      end

       2595 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2595");
      end

       2596 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2596");
      end

       2597 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2597");
      end

       2598 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2598");
      end

       2599 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2599");
      end

       2600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2600");
      end

       2601 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2601");
      end

       2602 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2602");
      end

       2603 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2603");
      end

       2604 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2604");
      end

       2605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2605");
      end

       2606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2606");
      end

       2607 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2607");
      end

       2608 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2608");
      end

       2609 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2609");
      end

       2610 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2610");
      end

       2611 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2611");
      end

       2612 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2612");
      end

       2613 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2613");
      end

       2614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2614");
      end

       2615 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2615");
      end

       2616 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2616");
      end

       2617 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2617");
      end

       2618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2618");
      end

       2619 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2619");
      end

       2620 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2620");
      end

       2621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2621");
      end

       2622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2622");
      end

       2623 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2623");
      end

       2624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2624");
      end

       2625 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2625");
      end

       2626 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2626");
      end

       2627 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2627");
      end

       2628 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2628");
      end

       2629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2629");
      end

       2630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2630");
      end

       2631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2631");
      end

       2632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2632");
      end

       2633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2633");
      end

       2634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2634");
      end

       2635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2635");
      end

       2636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2636");
      end

       2637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2637");
      end

       2638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2638");
      end

       2639 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2639");
      end

       2640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2640");
      end

       2641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2641");
      end

       2642 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2642");
      end

       2643 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2643");
      end

       2644 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2644");
      end

       2645 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2645");
      end

       2646 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2646");
      end

       2647 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2647");
      end

       2648 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2648");
      end

       2649 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2649");
      end

       2650 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2650");
      end

       2651 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2651");
      end

       2652 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2652");
      end

       2653 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2653");
      end

       2654 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2654");
      end

       2655 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2655");
      end

       2656 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2656");
      end

       2657 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2657");
      end

       2658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2658");
      end

       2659 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2659");
      end

       2660 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2660");
      end

       2661 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2661");
      end

       2662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2662");
      end

       2663 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  2663");
      end

       2664 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2664");
      end

       2665 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2665");
      end

       2666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2666");
      end

       2667 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2667");
      end

       2668 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2668");
      end

       2669 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2669");
      end

       2670 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  2670");
      end

       2671 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2671");
      end

       2672 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2672");
      end

       2673 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2673");
      end

       2674 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2674");
      end

       2675 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2675");
      end

       2676 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2676");
      end

       2677 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2677");
      end

       2678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2678");
      end

       2679 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2679");
      end

       2680 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2680");
      end

       2681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2681");
      end

       2682 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2682");
      end

       2683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2683");
      end

       2684 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  2684");
      end

       2685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2685");
      end

       2686 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  2686");
      end

       2687 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2687");
      end

       2688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2688");
      end

       2689 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2689");
      end

       2690 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2690");
      end

       2691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2691");
      end

       2692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2692");
      end

       2693 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2693");
      end

       2694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2694");
      end

       2695 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2695");
      end

       2696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2696");
      end

       2697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2697");
      end

       2698 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2698");
      end

       2699 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2699");
      end

       2700 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2700");
      end

       2701 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2701");
      end

       2702 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2702");
      end

       2703 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2703");
      end

       2704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2704");
      end

       2705 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2705");
      end

       2706 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2706");
      end

       2707 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2707");
      end

       2708 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2708");
      end

       2709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2709");
      end

       2710 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2710");
      end

       2711 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2711");
      end

       2712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2712");
      end

       2713 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2713");
      end

       2714 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2714");
      end

       2715 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2715");
      end

       2716 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2716");
      end

       2717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2717");
      end

       2718 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2718");
      end

       2719 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2719");
      end

       2720 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2720");
      end

       2721 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2721");
      end

       2722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2722");
      end

       2723 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2723");
      end

       2724 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2724");
      end

       2725 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2725");
      end

       2726 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2726");
      end

       2727 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2727");
      end

       2728 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2728");
      end

       2729 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2729");
      end

       2730 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2730");
      end

       2731 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2731");
      end

       2732 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2732");
      end

       2733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2733");
      end

       2734 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2734");
      end

       2735 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2735");
      end

       2736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2736");
      end

       2737 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2737");
      end

       2738 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2738");
      end

       2739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2739");
      end

       2740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2740");
      end

       2741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2741");
      end

       2742 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2742");
      end

       2743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2743");
      end

       2744 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2744");
      end

       2745 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2745");
      end

       2746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2746");
      end

       2747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2747");
      end

       2748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2748");
      end

       2749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2749");
      end

       2750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2750");
      end

       2751 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2751");
      end

       2752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2752");
      end

       2753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2753");
      end

       2754 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2754");
      end

       2755 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2755");
      end

       2756 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2756");
      end

       2757 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2757");
      end

       2758 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2758");
      end

       2759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2759");
      end

       2760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2760");
      end

       2761 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2761");
      end

       2762 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2762");
      end

       2763 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2763");
      end

       2764 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  2764");
      end

       2765 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2765");
      end

       2766 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  2766");
      end

       2767 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  2767");
      end

       2768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2768");
      end

       2769 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2769");
      end

       2770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2770");
      end

       2771 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2771");
      end

       2772 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2772");
      end

       2773 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2773");
      end

       2774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2774");
      end

       2775 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2775");
      end

       2776 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2776");
      end

       2777 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2777");
      end

       2778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2778");
      end

       2779 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2779");
      end

       2780 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2780");
      end

       2781 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2781");
      end

       2782 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2782");
      end

       2783 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2783");
      end

       2784 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2784");
      end

       2785 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2785");
      end

       2786 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2786");
      end

       2787 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2787");
      end

       2788 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2788");
      end

       2789 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2789");
      end

       2790 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2790");
      end

       2791 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2791");
      end

       2792 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2792");
      end

       2793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2793");
      end

       2794 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2794");
      end

       2795 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2795");
      end

       2796 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2796");
      end

       2797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2797");
      end

       2798 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2798");
      end

       2799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2799");
      end

       2800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2800");
      end

       2801 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2801");
      end

       2802 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2802");
      end

       2803 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2803");
      end

       2804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2804");
      end

       2805 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2805");
      end

       2806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2806");
      end

       2807 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2807");
      end

       2808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2808");
      end

       2809 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2809");
      end

       2810 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2810");
      end

       2811 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2811");
      end

       2812 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2812");
      end

       2813 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2813");
      end

       2814 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2814");
      end

       2815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2815");
      end

       2816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2816");
      end

       2817 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2817");
      end

       2818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2818");
      end

       2819 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2819");
      end

       2820 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2820");
      end

       2821 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2821");
      end

       2822 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2822");
      end

       2823 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2823");
      end

       2824 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2824");
      end

       2825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2825");
      end

       2826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2826");
      end

       2827 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2827");
      end

       2828 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2828");
      end

       2829 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2829");
      end

       2830 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2830");
      end

       2831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2831");
      end

       2832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2832");
      end

       2833 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2833");
      end

       2834 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2834");
      end

       2835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2835");
      end

       2836 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2836");
      end

       2837 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2837");
      end

       2838 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2838");
      end

       2839 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2839");
      end

       2840 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2840");
      end

       2841 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2841");
      end

       2842 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2842");
      end

       2843 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2843");
      end

       2844 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2844");
      end

       2845 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2845");
      end

       2846 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2846");
      end

       2847 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2847");
      end

       2848 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2848");
      end

       2849 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2849");
      end

       2850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2850");
      end

       2851 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2851");
      end

       2852 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2852");
      end

       2853 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2853");
      end

       2854 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2854");
      end

       2855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2855");
      end

       2856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2856");
      end

       2857 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2857");
      end

       2858 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2858");
      end

       2859 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2859");
      end

       2860 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2860");
      end

       2861 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2861");
      end

       2862 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2862");
      end

       2863 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2863");
      end

       2864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2864");
      end

       2865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2865");
      end

       2866 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2866");
      end

       2867 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2867");
      end

       2868 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2868");
      end

       2869 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2869");
      end

       2870 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2870");
      end

       2871 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2871");
      end

       2872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2872");
      end

       2873 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2873");
      end

       2874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2874");
      end

       2875 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2875");
      end

       2876 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2876");
      end

       2877 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2877");
      end

       2878 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2878");
      end

       2879 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2879");
      end

       2880 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2880");
      end

       2881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2881");
      end

       2882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2882");
      end

       2883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2883");
      end

       2884 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2884");
      end

       2885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2885");
      end

       2886 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2886");
      end

       2887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2887");
      end

       2888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2888");
      end

       2889 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2889");
      end

       2890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2890");
      end

       2891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2891");
      end

       2892 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2892");
      end

       2893 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2893");
      end

       2894 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2894");
      end

       2895 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2895");
      end

       2896 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2896");
      end

       2897 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2897");
      end

       2898 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2898");
      end

       2899 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2899");
      end

       2900 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2900");
      end

       2901 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2901");
      end

       2902 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2902");
      end

       2903 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2903");
      end

       2904 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2904");
      end

       2905 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2905");
      end

       2906 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2906");
      end

       2907 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2907");
      end

       2908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2908");
      end

       2909 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2909");
      end

       2910 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2910");
      end

       2911 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2911");
      end

       2912 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2912");
      end

       2913 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2913");
      end

       2914 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
         $display("Should not be executed  2914");
      end

       2915 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2915");
      end

       2916 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2916");
      end

       2917 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2917");
      end

       2918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2918");
      end

       2919 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2919");
      end

       2920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2920");
      end

       2921 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2921");
      end

       2922 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2922");
      end

       2923 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2923");
      end

       2924 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2924");
      end

       2925 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2925");
      end

       2926 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2926");
      end

       2927 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2927");
      end

       2928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2928");
      end

       2929 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2929");
      end

       2930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2930");
      end

       2931 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2931");
      end

       2932 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2932");
      end

       2933 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2933");
      end

       2934 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2934");
      end

       2935 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2935");
      end

       2936 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2936");
      end

       2937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2937");
      end

       2938 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  2938");
      end

       2939 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2939");
      end

       2940 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2940");
      end

       2941 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2941");
      end

       2942 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2942");
      end

       2943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2943");
      end

       2944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2944");
      end

       2945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2945");
      end

       2946 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  2946");
      end

       2947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2947");
      end

       2948 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  2948");
      end

       2949 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2949");
      end

       2950 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2950");
      end

       2951 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  2951");
      end

       2952 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2952");
      end

       2953 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2953");
      end

       2954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2954");
      end

       2955 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2955");
      end

       2956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2956");
      end

       2957 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2957");
      end

       2958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2958");
      end

       2959 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2959");
      end

       2960 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2960");
      end

       2961 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2961");
      end

       2962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2962");
      end

       2963 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  2963");
      end

       2964 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  2964");
      end

       2965 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  2965");
      end

       2966 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2966");
      end

       2967 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2967");
      end

       2968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2968");
      end

       2969 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2969");
      end

       2970 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2970");
      end

       2971 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2971");
      end

       2972 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2972");
      end

       2973 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2973");
      end

       2974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2974");
      end

       2975 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2975");
      end

       2976 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2976");
      end

       2977 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2977");
      end

       2978 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2978");
      end

       2979 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2979");
      end

       2980 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2980");
      end

       2981 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2981");
      end

       2982 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2982");
      end

       2983 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  2983");
      end

       2984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2984");
      end

       2985 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2985");
      end

       2986 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2986");
      end

       2987 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  2987");
      end

       2988 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2988");
      end

       2989 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2989");
      end

       2990 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2990");
      end

       2991 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  2991");
      end

       2992 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  2992");
      end

       2993 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  2993");
      end

       2994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2994");
      end

       2995 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2995");
      end

       2996 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2996");
      end

       2997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2997");
      end

       2998 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  2998");
      end

       2999 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  2999");
      end

       3000 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3000");
      end

       3001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3001");
      end

       3002 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3002");
      end

       3003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3003");
      end

       3004 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3004");
      end

       3005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3005");
      end

       3006 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3006");
      end

       3007 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3007");
      end

       3008 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3008");
      end

       3009 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3009");
      end

       3010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3010");
      end

       3011 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3011");
      end

       3012 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3012");
      end

       3013 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3013");
      end

       3014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3014");
      end

       3015 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3015");
      end

       3016 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3016");
      end

       3017 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3017");
      end

       3018 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3018");
      end

       3019 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3019");
      end

       3020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3020");
      end

       3021 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3021");
      end

       3022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3022");
      end

       3023 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3023");
      end

       3024 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3024");
      end

       3025 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3025");
      end

       3026 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  3026");
      end

       3027 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3027");
      end

       3028 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  3028");
      end

       3029 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  3029");
      end

       3030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3030");
      end

       3031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3031");
      end

       3032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3032");
      end

       3033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3033");
      end

       3034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3034");
      end

       3035 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3035");
      end

       3036 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3036");
      end

       3037 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3037");
      end

       3038 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3038");
      end

       3039 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3039");
      end

       3040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3040");
      end

       3041 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3041");
      end

       3042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3042");
      end

       3043 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3043");
      end

       3044 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3044");
      end

       3045 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3045");
      end

       3046 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3046");
      end

       3047 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3047");
      end

       3048 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3048");
      end

       3049 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3049");
      end

       3050 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3050");
      end

       3051 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3051");
      end

       3052 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3052");
      end

       3053 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3053");
      end

       3054 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3054");
      end

       3055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3055");
      end

       3056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3056");
      end

       3057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3057");
      end

       3058 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3058");
      end

       3059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3059");
      end

       3060 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3060");
      end

       3061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3061");
      end

       3062 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3062");
      end

       3063 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3063");
      end

       3064 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3064");
      end

       3065 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3065");
      end

       3066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3066");
      end

       3067 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3067");
      end

       3068 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3068");
      end

       3069 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3069");
      end

       3070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3070");
      end

       3071 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3071");
      end

       3072 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3072");
      end

       3073 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3073");
      end

       3074 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3074");
      end

       3075 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3075");
      end

       3076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3076");
      end

       3077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3077");
      end

       3078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3078");
      end

       3079 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3079");
      end

       3080 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3080");
      end

       3081 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3081");
      end

       3082 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3082");
      end

       3083 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3083");
      end

       3084 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3084");
      end

       3085 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3085");
      end

       3086 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3086");
      end

       3087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3087");
      end

       3088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3088");
      end

       3089 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3089");
      end

       3090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3090");
      end

       3091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3091");
      end

       3092 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3092");
      end

       3093 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3093");
      end

       3094 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3094");
      end

       3095 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3095");
      end

       3096 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3096");
      end

       3097 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3097");
      end

       3098 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3098");
      end

       3099 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3099");
      end

       3100 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3100");
      end

       3101 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3101");
      end

       3102 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3102");
      end

       3103 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3103");
      end

       3104 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3104");
      end

       3105 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3105");
      end

       3106 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3106");
      end

       3107 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3107");
      end

       3108 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3108");
      end

       3109 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3109");
      end

       3110 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3110");
      end

       3111 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3111");
      end

       3112 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3112");
      end

       3113 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3113");
      end

       3114 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3114");
      end

       3115 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3115");
      end

       3116 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3116");
      end

       3117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3117");
      end

       3118 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3118");
      end

       3119 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3119");
      end

       3120 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3120");
      end

       3121 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3121");
      end

       3122 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3122");
      end

       3123 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3123");
      end

       3124 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3124");
      end

       3125 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3125");
      end

       3126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3126");
      end

       3127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3127");
      end

       3128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3128");
      end

       3129 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3129");
      end

       3130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3130");
      end

       3131 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3131");
      end

       3132 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3132");
      end

       3133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3133");
      end

       3134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3134");
      end

       3135 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3135");
      end

       3136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3136");
      end

       3137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3137");
      end

       3138 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3138");
      end

       3139 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3139");
      end

       3140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3140");
      end

       3141 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3141");
      end

       3142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3142");
      end

       3143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3143");
      end

       3144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3144");
      end

       3145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3145");
      end

       3146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3146");
      end

       3147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3147");
      end

       3148 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3148");
      end

       3149 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3149");
      end

       3150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3150");
      end

       3151 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3151");
      end

       3152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3152");
      end

       3153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3153");
      end

       3154 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3154");
      end

       3155 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3155");
      end

       3156 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3156");
      end

       3157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3157");
      end

       3158 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3158");
      end

       3159 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3159");
      end

       3160 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3160");
      end

       3161 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3161");
      end

       3162 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3162");
      end

       3163 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3163");
      end

       3164 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3164");
      end

       3165 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3165");
      end

       3166 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3166");
      end

       3167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3167");
      end

       3168 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3168");
      end

       3169 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3169");
      end

       3170 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3170");
      end

       3171 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3172;
      end

       3172 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[951]] = 0;
              freedArrays[freedArraysTop] = localMem[951];
              freedArraysTop = freedArraysTop + 1;
              ip = 3173;
      end

       3173 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1426] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1426] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1426]] = 0;
              ip = 3174;
      end

       3174 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3175;
      end

       3175 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1427] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3176;
      end

       3176 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1427] != 0 ? 3199 : 3177;
      end

       3177 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3177");
      end

       3178 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3178");
      end

       3179 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3179");
      end

       3180 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3180");
      end

       3181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3181");
      end

       3182 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3182");
      end

       3183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3183");
      end

       3184 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3184");
      end

       3185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3185");
      end

       3186 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3186");
      end

       3187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3187");
      end

       3188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3188");
      end

       3189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3189");
      end

       3190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3190");
      end

       3191 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3191");
      end

       3192 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3192");
      end

       3193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3193");
      end

       3194 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3194");
      end

       3195 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3195");
      end

       3196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3196");
      end

       3197 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3197");
      end

       3198 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3198");
      end

       3199 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3200;
      end

       3200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1435] = heapMem[localMem[1427]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3201;
      end

       3201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1436] = heapMem[localMem[0]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3202;
      end

       3202 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1435] >= localMem[1436] ? 3238 : 3203;
      end

       3203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3203");
      end

       3204 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3204");
      end

       3205 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3205");
      end

       3206 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  3206");
      end

       3207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3207");
      end

       3208 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  3208");
      end

       3209 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  3209");
      end

       3210 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  3210");
      end

       3211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3211");
      end

       3212 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3212");
      end

       3213 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3213");
      end

       3214 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3214");
      end

       3215 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3215");
      end

       3216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3216");
      end

       3217 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3217");
      end

       3218 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
         $display("Should not be executed  3218");
      end

       3219 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3219");
      end

       3220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3220");
      end

       3221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3221");
      end

       3222 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3222");
      end

       3223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3223");
      end

       3224 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3224");
      end

       3225 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3225");
      end

       3226 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3226");
      end

       3227 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3227");
      end

       3228 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  3228");
      end

       3229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3229");
      end

       3230 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3230");
      end

       3231 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3231");
      end

       3232 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3232");
      end

       3233 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3233");
      end

       3234 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3234");
      end

       3235 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3235");
      end

       3236 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3236");
      end

       3237 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3237");
      end

       3238 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3239;
      end

       3239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1449] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3240;
      end

       3240 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3241;
      end

       3241 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1451] = heapMem[localMem[1449]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3242;
      end

       3242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1452] = heapMem[localMem[1449]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3243;
      end

       3243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1453] = heapMem[localMem[1452]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3244;
      end

       3244 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1451] <  localMem[1453] ? 3464 : 3245;
      end

       3245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1454] = localMem[1453];
              updateArrayLength(2, 0, 0);
              ip = 3246;
      end

       3246 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[1454] = localMem[1454] >> 1;
              ip = 3247;
      end

       3247 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1455] = localMem[1454] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3248;
      end

       3248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1456] = heapMem[localMem[1449]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3249;
      end

       3249 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1456] == 0 ? 3346 : 3250;
      end

       3250 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3250");
      end

       3251 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3251");
      end

       3252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3252");
      end

       3253 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3253");
      end

       3254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3254");
      end

       3255 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3255");
      end

       3256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3256");
      end

       3257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3257");
      end

       3258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3258");
      end

       3259 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3259");
      end

       3260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3260");
      end

       3261 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3261");
      end

       3262 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3262");
      end

       3263 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3263");
      end

       3264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3264");
      end

       3265 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3265");
      end

       3266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3266");
      end

       3267 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3267");
      end

       3268 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3268");
      end

       3269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3269");
      end

       3270 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3270");
      end

       3271 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3271");
      end

       3272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3272");
      end

       3273 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3273");
      end

       3274 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3274");
      end

       3275 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3275");
      end

       3276 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3276");
      end

       3277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3277");
      end

       3278 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3278");
      end

       3279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3279");
      end

       3280 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3280");
      end

       3281 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3281");
      end

       3282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3282");
      end

       3283 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3283");
      end

       3284 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3284");
      end

       3285 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3285");
      end

       3286 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3286");
      end

       3287 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3287");
      end

       3288 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3288");
      end

       3289 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3289");
      end

       3290 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3290");
      end

       3291 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3291");
      end

       3292 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3292");
      end

       3293 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3293");
      end

       3294 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3294");
      end

       3295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3295");
      end

       3296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3296");
      end

       3297 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3297");
      end

       3298 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3298");
      end

       3299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3299");
      end

       3300 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3300");
      end

       3301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3301");
      end

       3302 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3302");
      end

       3303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3303");
      end

       3304 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3304");
      end

       3305 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3305");
      end

       3306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3306");
      end

       3307 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3307");
      end

       3308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3308");
      end

       3309 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3309");
      end

       3310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3310");
      end

       3311 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3311");
      end

       3312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3312");
      end

       3313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3313");
      end

       3314 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3314");
      end

       3315 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3315");
      end

       3316 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3316");
      end

       3317 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3317");
      end

       3318 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3318");
      end

       3319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3319");
      end

       3320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3320");
      end

       3321 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3321");
      end

       3322 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3322");
      end

       3323 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3323");
      end

       3324 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  3324");
      end

       3325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3325");
      end

       3326 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  3326");
      end

       3327 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  3327");
      end

       3328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3328");
      end

       3329 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3329");
      end

       3330 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3330");
      end

       3331 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3331");
      end

       3332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3332");
      end

       3333 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3333");
      end

       3334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3334");
      end

       3335 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3335");
      end

       3336 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3336");
      end

       3337 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3337");
      end

       3338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3338");
      end

       3339 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3339");
      end

       3340 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3340");
      end

       3341 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3341");
      end

       3342 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3342");
      end

       3343 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3343");
      end

       3344 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3344");
      end

       3345 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3345");
      end

       3346 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3347;
      end

       3347 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1504] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1504] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1504]] = 0;
              ip = 3348;
      end

       3348 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 0] = localMem[1454];
              updateArrayLength(1, localMem[1504], 0);
              ip = 3349;
      end

       3349 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 2] = 0;
              updateArrayLength(1, localMem[1504], 2);
              ip = 3350;
      end

       3350 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1505] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1505] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1505]] = 0;
              ip = 3351;
      end

       3351 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 4] = localMem[1505];
              updateArrayLength(1, localMem[1504], 4);
              ip = 3352;
      end

       3352 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1506] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1506] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1506]] = 0;
              ip = 3353;
      end

       3353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 5] = localMem[1506];
              updateArrayLength(1, localMem[1504], 5);
              ip = 3354;
      end

       3354 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 6] = 0;
              updateArrayLength(1, localMem[1504], 6);
              ip = 3355;
      end

       3355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 3] = localMem[1452];
              updateArrayLength(1, localMem[1504], 3);
              ip = 3356;
      end

       3356 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1452]*7 + 1] = heapMem[localMem[1452]*7 + 1] + 1;
              updateArrayLength(1, localMem[1452], 1);
              ip = 3357;
      end

       3357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 1] = heapMem[localMem[1452]*7 + 1];
              updateArrayLength(1, localMem[1504], 1);
              ip = 3358;
      end

       3358 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1507] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1507] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1507]] = 0;
              ip = 3359;
      end

       3359 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 0] = localMem[1454];
              updateArrayLength(1, localMem[1507], 0);
              ip = 3360;
      end

       3360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 2] = 0;
              updateArrayLength(1, localMem[1507], 2);
              ip = 3361;
      end

       3361 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1508] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1508] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1508]] = 0;
              ip = 3362;
      end

       3362 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 4] = localMem[1508];
              updateArrayLength(1, localMem[1507], 4);
              ip = 3363;
      end

       3363 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1509] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1509] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1509]] = 0;
              ip = 3364;
      end

       3364 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 5] = localMem[1509];
              updateArrayLength(1, localMem[1507], 5);
              ip = 3365;
      end

       3365 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 6] = 0;
              updateArrayLength(1, localMem[1507], 6);
              ip = 3366;
      end

       3366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 3] = localMem[1452];
              updateArrayLength(1, localMem[1507], 3);
              ip = 3367;
      end

       3367 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1452]*7 + 1] = heapMem[localMem[1452]*7 + 1] + 1;
              updateArrayLength(1, localMem[1452], 1);
              ip = 3368;
      end

       3368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 1] = heapMem[localMem[1452]*7 + 1];
              updateArrayLength(1, localMem[1507], 1);
              ip = 3369;
      end

       3369 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1510] = !heapMem[localMem[1449]*7 + 6];
              ip = 3370;
      end

       3370 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1510] != 0 ? 3422 : 3371;
      end

       3371 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3371");
      end

       3372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3372");
      end

       3373 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3373");
      end

       3374 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3374");
      end

       3375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3375");
      end

       3376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3376");
      end

       3377 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3377");
      end

       3378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3378");
      end

       3379 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3379");
      end

       3380 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3380");
      end

       3381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3381");
      end

       3382 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3382");
      end

       3383 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3383");
      end

       3384 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3384");
      end

       3385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3385");
      end

       3386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3386");
      end

       3387 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3387");
      end

       3388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3388");
      end

       3389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3389");
      end

       3390 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3390");
      end

       3391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3391");
      end

       3392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3392");
      end

       3393 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3393");
      end

       3394 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3394");
      end

       3395 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3395");
      end

       3396 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3396");
      end

       3397 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3397");
      end

       3398 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3398");
      end

       3399 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3399");
      end

       3400 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3400");
      end

       3401 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3401");
      end

       3402 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3402");
      end

       3403 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3403");
      end

       3404 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3404");
      end

       3405 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3405");
      end

       3406 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3406");
      end

       3407 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3407");
      end

       3408 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3408");
      end

       3409 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3409");
      end

       3410 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3410");
      end

       3411 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3411");
      end

       3412 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3412");
      end

       3413 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3413");
      end

       3414 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3414");
      end

       3415 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3415");
      end

       3416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3416");
      end

       3417 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3417");
      end

       3418 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3418");
      end

       3419 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3419");
      end

       3420 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3420");
      end

       3421 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3421");
      end

       3422 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3423;
      end

       3423 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1537] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1537] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1537]] = 0;
              ip = 3424;
      end

       3424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1449]*7 + 6] = localMem[1537];
              updateArrayLength(1, localMem[1449], 6);
              ip = 3425;
      end

       3425 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1538] = heapMem[localMem[1449]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3426;
      end

       3426 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1539] = heapMem[localMem[1504]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3427;
      end

       3427 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1539] + 0 + i] = heapMem[NArea * localMem[1538] + 0 + i];
                  updateArrayLength(1, localMem[1539], 0 + i);
                end
              end
              ip = 3428;
      end

       3428 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1540] = heapMem[localMem[1449]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3429;
      end

       3429 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1541] = heapMem[localMem[1504]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3430;
      end

       3430 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1541] + 0 + i] = heapMem[NArea * localMem[1540] + 0 + i];
                  updateArrayLength(1, localMem[1541], 0 + i);
                end
              end
              ip = 3431;
      end

       3431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1542] = heapMem[localMem[1449]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3432;
      end

       3432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1543] = heapMem[localMem[1507]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3433;
      end

       3433 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1543] + 0 + i] = heapMem[NArea * localMem[1542] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1543], 0 + i);
                end
              end
              ip = 3434;
      end

       3434 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1544] = heapMem[localMem[1449]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3435;
      end

       3435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1545] = heapMem[localMem[1507]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3436;
      end

       3436 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[1454]) begin
                  heapMem[NArea * localMem[1545] + 0 + i] = heapMem[NArea * localMem[1544] + localMem[1455] + i];
                  updateArrayLength(1, localMem[1545], 0 + i);
                end
              end
              ip = 3437;
      end

       3437 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3438;
      end

       3438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1504]*7 + 2] = localMem[1449];
              updateArrayLength(1, localMem[1504], 2);
              ip = 3439;
      end

       3439 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1507]*7 + 2] = localMem[1449];
              updateArrayLength(1, localMem[1507], 2);
              ip = 3440;
      end

       3440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1546] = heapMem[localMem[1449]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3441;
      end

       3441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1547] = heapMem[localMem[1546]*7 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3442;
      end

       3442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1548] = heapMem[localMem[1449]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3443;
      end

       3443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1549] = heapMem[localMem[1548]*7 + localMem[1454]];
              updateArrayLength(2, 0, 0);
              ip = 3444;
      end

       3444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1550] = heapMem[localMem[1449]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3445;
      end

       3445 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1550]*7 + 0] = localMem[1547];
              updateArrayLength(1, localMem[1550], 0);
              ip = 3446;
      end

       3446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1551] = heapMem[localMem[1449]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3447;
      end

       3447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1551]*7 + 0] = localMem[1549];
              updateArrayLength(1, localMem[1551], 0);
              ip = 3448;
      end

       3448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1552] = heapMem[localMem[1449]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3449;
      end

       3449 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1552]*7 + 0] = localMem[1504];
              updateArrayLength(1, localMem[1552], 0);
              ip = 3450;
      end

       3450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1553] = heapMem[localMem[1449]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3451;
      end

       3451 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1553]*7 + 1] = localMem[1507];
              updateArrayLength(1, localMem[1553], 1);
              ip = 3452;
      end

       3452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1449]*7 + 0] = 1;
              updateArrayLength(1, localMem[1449], 0);
              ip = 3453;
      end

       3453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1554] = heapMem[localMem[1449]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3454;
      end

       3454 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1554]] = 1;
              ip = 3455;
      end

       3455 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1555] = heapMem[localMem[1449]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3456;
      end

       3456 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1555]] = 1;
              ip = 3457;
      end

       3457 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1556] = heapMem[localMem[1449]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3458;
      end

       3458 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[1556]] = 2;
              ip = 3459;
      end

       3459 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3461;
      end

       3460 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3460");
      end

       3461 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3462;
      end

       3462 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1450] = 1;
              updateArrayLength(2, 0, 0);
              ip = 3463;
      end

       3463 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3466;
      end

       3464 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3464");
      end

       3465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3465");
      end

       3466 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3467;
      end

       3467 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3468;
      end

       3468 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3469;
      end

       3469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1557] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3470;
      end

       3470 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3471;
      end

       3471 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1557] >= 99 ? 3969 : 3472;
      end

       3472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1558] = heapMem[localMem[1449]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3473;
      end

       3473 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[1559] = localMem[1558] - 1;
              updateArrayLength(2, 0, 0);
              ip = 3474;
      end

       3474 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1560] = heapMem[localMem[1449]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3475;
      end

       3475 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1561] = heapMem[localMem[1560]*7 + localMem[1559]];
              updateArrayLength(2, 0, 0);
              ip = 3476;
      end

       3476 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 4 <= localMem[1561] ? 3717 : 3477;
      end

       3477 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1562] = !heapMem[localMem[1449]*7 + 6];
              ip = 3478;
      end

       3478 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1562] == 0 ? 3483 : 3479;
      end

       3479 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*7 + 0] = localMem[1449];
              updateArrayLength(1, localMem[1426], 0);
              ip = 3480;
      end

       3480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1426]*7 + 1] = 2;
              updateArrayLength(1, localMem[1426], 1);
              ip = 3481;
      end

       3481 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1426]*7 + 2] = localMem[1558] - 1;
              updateArrayLength(1, localMem[1426], 2);
              ip = 3482;
      end

       3482 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3973;
      end

       3483 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3484;
      end

       3484 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1563] = heapMem[localMem[1449]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 3485;
      end

       3485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1564] = heapMem[localMem[1563]*7 + localMem[1558]];
              updateArrayLength(2, 0, 0);
              ip = 3486;
      end

       3486 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3487;
      end

       3487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1566] = heapMem[localMem[1564]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3488;
      end

       3488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1567] = heapMem[localMem[1564]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 3489;
      end

       3489 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1568] = heapMem[localMem[1567]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3490;
      end

       3490 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1566] <  localMem[1568] ? 3710 : 3491;
      end

       3491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3491");
      end

       3492 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  3492");
      end

       3493 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3493");
      end

       3494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3494");
      end

       3495 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  3495");
      end

       3496 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3496");
      end

       3497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3497");
      end

       3498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3498");
      end

       3499 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3499");
      end

       3500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3500");
      end

       3501 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3501");
      end

       3502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3502");
      end

       3503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3503");
      end

       3504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3504");
      end

       3505 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3505");
      end

       3506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3506");
      end

       3507 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3507");
      end

       3508 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3508");
      end

       3509 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3509");
      end

       3510 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3510");
      end

       3511 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3511");
      end

       3512 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3512");
      end

       3513 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3513");
      end

       3514 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3514");
      end

       3515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3515");
      end

       3516 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3516");
      end

       3517 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3517");
      end

       3518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3518");
      end

       3519 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3519");
      end

       3520 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3520");
      end

       3521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3521");
      end

       3522 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3522");
      end

       3523 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3523");
      end

       3524 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3524");
      end

       3525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3525");
      end

       3526 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3526");
      end

       3527 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3527");
      end

       3528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3528");
      end

       3529 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3529");
      end

       3530 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3530");
      end

       3531 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3531");
      end

       3532 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3532");
      end

       3533 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3533");
      end

       3534 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3534");
      end

       3535 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3535");
      end

       3536 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3536");
      end

       3537 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3537");
      end

       3538 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3538");
      end

       3539 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3539");
      end

       3540 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3540");
      end

       3541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3541");
      end

       3542 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3542");
      end

       3543 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3543");
      end

       3544 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3544");
      end

       3545 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3545");
      end

       3546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3546");
      end

       3547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3547");
      end

       3548 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3548");
      end

       3549 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3549");
      end

       3550 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3550");
      end

       3551 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3551");
      end

       3552 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3552");
      end

       3553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3553");
      end

       3554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3554");
      end

       3555 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3555");
      end

       3556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3556");
      end

       3557 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3557");
      end

       3558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3558");
      end

       3559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3559");
      end

       3560 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3560");
      end

       3561 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3561");
      end

       3562 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3562");
      end

       3563 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3563");
      end

       3564 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3564");
      end

       3565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3565");
      end

       3566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3566");
      end

       3567 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3567");
      end

       3568 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3568");
      end

       3569 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3569");
      end

       3570 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  3570");
      end

       3571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3571");
      end

       3572 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  3572");
      end

       3573 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  3573");
      end

       3574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3574");
      end

       3575 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3575");
      end

       3576 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3576");
      end

       3577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3577");
      end

       3578 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3578");
      end

       3579 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3579");
      end

       3580 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3580");
      end

       3581 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3581");
      end

       3582 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3582");
      end

       3583 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3583");
      end

       3584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3584");
      end

       3585 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3585");
      end

       3586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3586");
      end

       3587 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3587");
      end

       3588 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3588");
      end

       3589 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3589");
      end

       3590 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3590");
      end

       3591 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3591");
      end

       3592 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3592");
      end

       3593 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3593");
      end

       3594 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3594");
      end

       3595 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3595");
      end

       3596 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3596");
      end

       3597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3597");
      end

       3598 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3598");
      end

       3599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3599");
      end

       3600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3600");
      end

       3601 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3601");
      end

       3602 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3602");
      end

       3603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3603");
      end

       3604 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3604");
      end

       3605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3605");
      end

       3606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3606");
      end

       3607 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3607");
      end

       3608 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3608");
      end

       3609 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3609");
      end

       3610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3610");
      end

       3611 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3611");
      end

       3612 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3612");
      end

       3613 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3613");
      end

       3614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3614");
      end

       3615 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3615");
      end

       3616 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3616");
      end

       3617 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3617");
      end

       3618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3618");
      end

       3619 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3619");
      end

       3620 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3620");
      end

       3621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3621");
      end

       3622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3622");
      end

       3623 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3623");
      end

       3624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3624");
      end

       3625 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3625");
      end

       3626 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3626");
      end

       3627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3627");
      end

       3628 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3628");
      end

       3629 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3629");
      end

       3630 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3630");
      end

       3631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3631");
      end

       3632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3632");
      end

       3633 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3633");
      end

       3634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3634");
      end

       3635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3635");
      end

       3636 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3636");
      end

       3637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3637");
      end

       3638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3638");
      end

       3639 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3639");
      end

       3640 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3640");
      end

       3641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3641");
      end

       3642 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3642");
      end

       3643 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3643");
      end

       3644 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3644");
      end

       3645 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3645");
      end

       3646 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3646");
      end

       3647 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3647");
      end

       3648 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3648");
      end

       3649 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3649");
      end

       3650 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3650");
      end

       3651 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3651");
      end

       3652 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3652");
      end

       3653 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3653");
      end

       3654 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3654");
      end

       3655 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3655");
      end

       3656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3656");
      end

       3657 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3657");
      end

       3658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3658");
      end

       3659 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3659");
      end

       3660 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3660");
      end

       3661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3661");
      end

       3662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3662");
      end

       3663 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3663");
      end

       3664 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3664");
      end

       3665 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3665");
      end

       3666 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3666");
      end

       3667 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3667");
      end

       3668 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3668");
      end

       3669 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3669");
      end

       3670 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3670");
      end

       3671 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3671");
      end

       3672 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3672");
      end

       3673 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3673");
      end

       3674 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3674");
      end

       3675 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3675");
      end

       3676 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3676");
      end

       3677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3677");
      end

       3678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3678");
      end

       3679 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3679");
      end

       3680 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3680");
      end

       3681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3681");
      end

       3682 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3682");
      end

       3683 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3683");
      end

       3684 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3684");
      end

       3685 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3685");
      end

       3686 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3686");
      end

       3687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3687");
      end

       3688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3688");
      end

       3689 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3689");
      end

       3690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3690");
      end

       3691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3691");
      end

       3692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3692");
      end

       3693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3693");
      end

       3694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3694");
      end

       3695 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3695");
      end

       3696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3696");
      end

       3697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3697");
      end

       3698 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3698");
      end

       3699 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3699");
      end

       3700 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3700");
      end

       3701 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3701");
      end

       3702 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3702");
      end

       3703 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3703");
      end

       3704 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3704");
      end

       3705 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3705");
      end

       3706 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3706");
      end

       3707 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3707");
      end

       3708 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3708");
      end

       3709 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3709");
      end

       3710 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3711;
      end

       3711 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1565] = 0;
              updateArrayLength(2, 0, 0);
              ip = 3712;
      end

       3712 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3713;
      end

       3713 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1565] != 0 ? 3715 : 3714;
      end

       3714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1449] = localMem[1564];
              updateArrayLength(2, 0, 0);
              ip = 3715;
      end

       3715 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3716;
      end

       3716 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3966;
      end

       3717 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3717");
      end

       3718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3718");
      end

       3719 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  3719");
      end

       3720 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  3720");
      end

       3721 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3721");
      end

       3722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3722");
      end

       3723 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  3723");
      end

       3724 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3724");
      end

       3725 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3725");
      end

       3726 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  3726");
      end

       3727 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3727");
      end

       3728 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  3728");
      end

       3729 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3729");
      end

       3730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3730");
      end

       3731 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3731");
      end

       3732 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3732");
      end

       3733 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3733");
      end

       3734 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3734");
      end

       3735 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3735");
      end

       3736 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3736");
      end

       3737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3737");
      end

       3738 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3738");
      end

       3739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3739");
      end

       3740 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  3740");
      end

       3741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3741");
      end

       3742 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  3742");
      end

       3743 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3743");
      end

       3744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3744");
      end

       3745 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  3745");
      end

       3746 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3746");
      end

       3747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3747");
      end

       3748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3748");
      end

       3749 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3749");
      end

       3750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3750");
      end

       3751 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3751");
      end

       3752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3752");
      end

       3753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3753");
      end

       3754 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3754");
      end

       3755 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3755");
      end

       3756 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3756");
      end

       3757 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3757");
      end

       3758 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3758");
      end

       3759 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3759");
      end

       3760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3760");
      end

       3761 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3761");
      end

       3762 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3762");
      end

       3763 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3763");
      end

       3764 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3764");
      end

       3765 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3765");
      end

       3766 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3766");
      end

       3767 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3767");
      end

       3768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3768");
      end

       3769 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3769");
      end

       3770 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3770");
      end

       3771 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3771");
      end

       3772 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3772");
      end

       3773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3773");
      end

       3774 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3774");
      end

       3775 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3775");
      end

       3776 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3776");
      end

       3777 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3777");
      end

       3778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3778");
      end

       3779 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3779");
      end

       3780 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3780");
      end

       3781 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3781");
      end

       3782 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3782");
      end

       3783 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3783");
      end

       3784 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3784");
      end

       3785 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3785");
      end

       3786 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3786");
      end

       3787 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3787");
      end

       3788 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3788");
      end

       3789 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3789");
      end

       3790 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3790");
      end

       3791 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3791");
      end

       3792 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3792");
      end

       3793 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3793");
      end

       3794 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3794");
      end

       3795 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3795");
      end

       3796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3796");
      end

       3797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3797");
      end

       3798 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3798");
      end

       3799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3799");
      end

       3800 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3800");
      end

       3801 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3801");
      end

       3802 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3802");
      end

       3803 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3803");
      end

       3804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3804");
      end

       3805 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3805");
      end

       3806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3806");
      end

       3807 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3807");
      end

       3808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3808");
      end

       3809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3809");
      end

       3810 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3810");
      end

       3811 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3811");
      end

       3812 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3812");
      end

       3813 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3813");
      end

       3814 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3814");
      end

       3815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3815");
      end

       3816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3816");
      end

       3817 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3817");
      end

       3818 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3818");
      end

       3819 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3819");
      end

       3820 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  3820");
      end

       3821 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3821");
      end

       3822 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  3822");
      end

       3823 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  3823");
      end

       3824 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3824");
      end

       3825 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3825");
      end

       3826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3826");
      end

       3827 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3827");
      end

       3828 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3828");
      end

       3829 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3829");
      end

       3830 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3830");
      end

       3831 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3831");
      end

       3832 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3832");
      end

       3833 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3833");
      end

       3834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3834");
      end

       3835 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3835");
      end

       3836 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3836");
      end

       3837 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3837");
      end

       3838 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3838");
      end

       3839 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3839");
      end

       3840 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3840");
      end

       3841 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3841");
      end

       3842 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3842");
      end

       3843 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3843");
      end

       3844 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3844");
      end

       3845 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3845");
      end

       3846 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3846");
      end

       3847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3847");
      end

       3848 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3848");
      end

       3849 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3849");
      end

       3850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3850");
      end

       3851 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3851");
      end

       3852 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3852");
      end

       3853 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3853");
      end

       3854 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3854");
      end

       3855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3855");
      end

       3856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3856");
      end

       3857 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3857");
      end

       3858 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3858");
      end

       3859 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3859");
      end

       3860 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3860");
      end

       3861 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3861");
      end

       3862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3862");
      end

       3863 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3863");
      end

       3864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3864");
      end

       3865 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  3865");
      end

       3866 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3866");
      end

       3867 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3867");
      end

       3868 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3868");
      end

       3869 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3869");
      end

       3870 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3870");
      end

       3871 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3871");
      end

       3872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3872");
      end

       3873 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3873");
      end

       3874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3874");
      end

       3875 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3875");
      end

       3876 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3876");
      end

       3877 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3877");
      end

       3878 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3878");
      end

       3879 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3879");
      end

       3880 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3880");
      end

       3881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3881");
      end

       3882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3882");
      end

       3883 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3883");
      end

       3884 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3884");
      end

       3885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3885");
      end

       3886 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3886");
      end

       3887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3887");
      end

       3888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3888");
      end

       3889 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3889");
      end

       3890 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3890");
      end

       3891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3891");
      end

       3892 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3892");
      end

       3893 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3893");
      end

       3894 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3894");
      end

       3895 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3895");
      end

       3896 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3896");
      end

       3897 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3897");
      end

       3898 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3898");
      end

       3899 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3899");
      end

       3900 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3900");
      end

       3901 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3901");
      end

       3902 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3902");
      end

       3903 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3903");
      end

       3904 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3904");
      end

       3905 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3905");
      end

       3906 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3906");
      end

       3907 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3907");
      end

       3908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3908");
      end

       3909 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3909");
      end

       3910 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  3910");
      end

       3911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3911");
      end

       3912 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3912");
      end

       3913 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3913");
      end

       3914 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3914");
      end

       3915 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3915");
      end

       3916 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3916");
      end

       3917 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3917");
      end

       3918 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3918");
      end

       3919 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  3919");
      end

       3920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3920");
      end

       3921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3921");
      end

       3922 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3922");
      end

       3923 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3923");
      end

       3924 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3924");
      end

       3925 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3925");
      end

       3926 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3926");
      end

       3927 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3927");
      end

       3928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3928");
      end

       3929 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3929");
      end

       3930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3930");
      end

       3931 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3931");
      end

       3932 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  3932");
      end

       3933 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3933");
      end

       3934 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3934");
      end

       3935 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3935");
      end

       3936 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3936");
      end

       3937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3937");
      end

       3938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3938");
      end

       3939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3939");
      end

       3940 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3940");
      end

       3941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3941");
      end

       3942 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3942");
      end

       3943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3943");
      end

       3944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3944");
      end

       3945 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3945");
      end

       3946 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3946");
      end

       3947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3947");
      end

       3948 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3948");
      end

       3949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3949");
      end

       3950 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3950");
      end

       3951 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3951");
      end

       3952 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3952");
      end

       3953 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3953");
      end

       3954 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  3954");
      end

       3955 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3955");
      end

       3956 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3956");
      end

       3957 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3957");
      end

       3958 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3958");
      end

       3959 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3959");
      end

       3960 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3960");
      end

       3961 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3961");
      end

       3962 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3962");
      end

       3963 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  3963");
      end

       3964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3964");
      end

       3965 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3965");
      end

       3966 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3967;
      end

       3967 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1557] = localMem[1557] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3968;
      end

       3968 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3470;
      end

       3969 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3969");
      end

       3970 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
         $display("Should not be executed  3970");
      end

       3971 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3971");
      end

       3972 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3972");
      end

       3973 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3974;
      end

       3974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1785] = heapMem[localMem[1426]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 3975;
      end

       3975 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1786] = heapMem[localMem[1426]*7 + 1];
              updateArrayLength(2, 0, 0);
              ip = 3976;
      end

       3976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1787] = heapMem[localMem[1426]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 3977;
      end

       3977 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1786] != 1 ? 3981 : 3978;
      end

       3978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3978");
      end

       3979 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3979");
      end

       3980 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  3980");
      end

       3981 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3982;
      end

       3982 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1786] != 2 ? 3990 : 3983;
      end

       3983 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[1789] = localMem[1787] + 1;
              updateArrayLength(2, 0, 0);
              ip = 3984;
      end

       3984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1790] = heapMem[localMem[1785]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 3985;
      end

       3985 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1790] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1789], localMem[1790], arraySizes[localMem[1790]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1789] && i <= arraySizes[localMem[1790]]) begin
                  heapMem[NArea * localMem[1790] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1790] + localMem[1789]] = 4;                                    // Insert new value
              arraySizes[localMem[1790]] = arraySizes[localMem[1790]] + 1;                              // Increase array size
              ip = 3986;
      end

       3986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1791] = heapMem[localMem[1785]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 3987;
      end

       3987 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[1791] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[1789], localMem[1791], arraySizes[localMem[1791]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[1789] && i <= arraySizes[localMem[1791]]) begin
                  heapMem[NArea * localMem[1791] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[1791] + localMem[1789]] = 44;                                    // Insert new value
              arraySizes[localMem[1791]] = arraySizes[localMem[1791]] + 1;                              // Increase array size
              ip = 3988;
      end

       3988 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[1785]*7 + 0] = heapMem[localMem[1785]*7 + 0] + 1;
              updateArrayLength(1, localMem[1785], 0);
              ip = 3989;
      end

       3989 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 3996;
      end

       3990 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  3990");
      end

       3991 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3991");
      end

       3992 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3992");
      end

       3993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  3993");
      end

       3994 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  3994");
      end

       3995 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  3995");
      end

       3996 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3997;
      end

       3997 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = heapMem[localMem[0]*7 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 3998;
      end

       3998 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 3999;
      end

       3999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1795] = heapMem[localMem[1785]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4000;
      end

       4000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1796] = heapMem[localMem[1785]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4001;
      end

       4001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1797] = heapMem[localMem[1796]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4002;
      end

       4002 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1795] <  localMem[1797] ? 4222 : 4003;
      end

       4003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4003");
      end

       4004 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  4004");
      end

       4005 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4005");
      end

       4006 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4006");
      end

       4007 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4007");
      end

       4008 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4008");
      end

       4009 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4009");
      end

       4010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4010");
      end

       4011 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4011");
      end

       4012 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4012");
      end

       4013 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4013");
      end

       4014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4014");
      end

       4015 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4015");
      end

       4016 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4016");
      end

       4017 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4017");
      end

       4018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4018");
      end

       4019 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4019");
      end

       4020 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4020");
      end

       4021 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4021");
      end

       4022 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4022");
      end

       4023 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4023");
      end

       4024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4024");
      end

       4025 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4025");
      end

       4026 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4026");
      end

       4027 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4027");
      end

       4028 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4028");
      end

       4029 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4029");
      end

       4030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4030");
      end

       4031 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4031");
      end

       4032 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4032");
      end

       4033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4033");
      end

       4034 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4034");
      end

       4035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4035");
      end

       4036 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4036");
      end

       4037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4037");
      end

       4038 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4038");
      end

       4039 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4039");
      end

       4040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4040");
      end

       4041 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4041");
      end

       4042 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4042");
      end

       4043 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4043");
      end

       4044 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4044");
      end

       4045 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4045");
      end

       4046 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4046");
      end

       4047 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4047");
      end

       4048 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4048");
      end

       4049 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4049");
      end

       4050 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4050");
      end

       4051 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4051");
      end

       4052 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4052");
      end

       4053 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4053");
      end

       4054 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4054");
      end

       4055 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4055");
      end

       4056 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4056");
      end

       4057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4057");
      end

       4058 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4058");
      end

       4059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4059");
      end

       4060 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4060");
      end

       4061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4061");
      end

       4062 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4062");
      end

       4063 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4063");
      end

       4064 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4064");
      end

       4065 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4065");
      end

       4066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4066");
      end

       4067 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4067");
      end

       4068 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4068");
      end

       4069 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4069");
      end

       4070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4070");
      end

       4071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4071");
      end

       4072 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4072");
      end

       4073 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4073");
      end

       4074 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4074");
      end

       4075 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4075");
      end

       4076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4076");
      end

       4077 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4077");
      end

       4078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4078");
      end

       4079 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4079");
      end

       4080 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4080");
      end

       4081 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4081");
      end

       4082 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  4082");
      end

       4083 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4083");
      end

       4084 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  4084");
      end

       4085 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  4085");
      end

       4086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4086");
      end

       4087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4087");
      end

       4088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4088");
      end

       4089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4089");
      end

       4090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4090");
      end

       4091 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4091");
      end

       4092 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4092");
      end

       4093 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4093");
      end

       4094 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4094");
      end

       4095 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4095");
      end

       4096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4096");
      end

       4097 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4097");
      end

       4098 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4098");
      end

       4099 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4099");
      end

       4100 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4100");
      end

       4101 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4101");
      end

       4102 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4102");
      end

       4103 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4103");
      end

       4104 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4104");
      end

       4105 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4105");
      end

       4106 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4106");
      end

       4107 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4107");
      end

       4108 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4108");
      end

       4109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4109");
      end

       4110 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4110");
      end

       4111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4111");
      end

       4112 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4112");
      end

       4113 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4113");
      end

       4114 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4114");
      end

       4115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4115");
      end

       4116 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4116");
      end

       4117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4117");
      end

       4118 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4118");
      end

       4119 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4119");
      end

       4120 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4120");
      end

       4121 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4121");
      end

       4122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4122");
      end

       4123 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4123");
      end

       4124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4124");
      end

       4125 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4125");
      end

       4126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4126");
      end

       4127 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4127");
      end

       4128 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4128");
      end

       4129 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4129");
      end

       4130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4130");
      end

       4131 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4131");
      end

       4132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4132");
      end

       4133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4133");
      end

       4134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4134");
      end

       4135 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4135");
      end

       4136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4136");
      end

       4137 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4137");
      end

       4138 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4138");
      end

       4139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4139");
      end

       4140 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4140");
      end

       4141 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4141");
      end

       4142 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4142");
      end

       4143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4143");
      end

       4144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4144");
      end

       4145 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4145");
      end

       4146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4146");
      end

       4147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4147");
      end

       4148 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4148");
      end

       4149 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4149");
      end

       4150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4150");
      end

       4151 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4151");
      end

       4152 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4152");
      end

       4153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4153");
      end

       4154 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4154");
      end

       4155 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4155");
      end

       4156 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4156");
      end

       4157 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4157");
      end

       4158 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4158");
      end

       4159 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4159");
      end

       4160 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4160");
      end

       4161 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4161");
      end

       4162 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4162");
      end

       4163 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4163");
      end

       4164 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4164");
      end

       4165 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4165");
      end

       4166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4166");
      end

       4167 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4167");
      end

       4168 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4168");
      end

       4169 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4169");
      end

       4170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4170");
      end

       4171 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4171");
      end

       4172 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4172");
      end

       4173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4173");
      end

       4174 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4174");
      end

       4175 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4175");
      end

       4176 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4176");
      end

       4177 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4177");
      end

       4178 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4178");
      end

       4179 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4179");
      end

       4180 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4180");
      end

       4181 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4181");
      end

       4182 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4182");
      end

       4183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4183");
      end

       4184 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4184");
      end

       4185 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4185");
      end

       4186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4186");
      end

       4187 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4187");
      end

       4188 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4188");
      end

       4189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4189");
      end

       4190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4190");
      end

       4191 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4191");
      end

       4192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4192");
      end

       4193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4193");
      end

       4194 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4194");
      end

       4195 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4195");
      end

       4196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4196");
      end

       4197 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4197");
      end

       4198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4198");
      end

       4199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4199");
      end

       4200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4200");
      end

       4201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4201");
      end

       4202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4202");
      end

       4203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4203");
      end

       4204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4204");
      end

       4205 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4205");
      end

       4206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4206");
      end

       4207 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4207");
      end

       4208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4208");
      end

       4209 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4209");
      end

       4210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4210");
      end

       4211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4211");
      end

       4212 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4212");
      end

       4213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4213");
      end

       4214 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4214");
      end

       4215 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4215");
      end

       4216 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4216");
      end

       4217 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4217");
      end

       4218 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4218");
      end

       4219 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4219");
      end

       4220 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4220");
      end

       4221 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4221");
      end

       4222 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4223;
      end

       4223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1794] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4224;
      end

       4224 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4225;
      end

       4225 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4226;
      end

       4226 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4227;
      end

       4227 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4228;
      end

       4228 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[1426]] = 0;
              freedArrays[freedArraysTop] = localMem[1426];
              freedArraysTop = freedArraysTop + 1;
              ip = 4229;
      end

       4229 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[1901] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[1901] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[1901]] = 0;
              ip = 4230;
      end

       4230 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4231;
      end

       4231 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1902] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4232;
      end

       4232 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1902] != 0 ? 4255 : 4233;
      end

       4233 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4233");
      end

       4234 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4234");
      end

       4235 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4235");
      end

       4236 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4236");
      end

       4237 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4237");
      end

       4238 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4238");
      end

       4239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4239");
      end

       4240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4240");
      end

       4241 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4241");
      end

       4242 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4242");
      end

       4243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4243");
      end

       4244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4244");
      end

       4245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4245");
      end

       4246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4246");
      end

       4247 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4247");
      end

       4248 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4248");
      end

       4249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4249");
      end

       4250 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4250");
      end

       4251 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4251");
      end

       4252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4252");
      end

       4253 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4253");
      end

       4254 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4254");
      end

       4255 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4256;
      end

       4256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1910] = heapMem[localMem[1902]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4257;
      end

       4257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1911] = heapMem[localMem[0]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4258;
      end

       4258 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[1910] >= localMem[1911] ? 4294 : 4259;
      end

       4259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1912] = heapMem[localMem[1902]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4260;
      end

       4260 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[1912] != 0 ? 4293 : 4261;
      end

       4261 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[1913] = !heapMem[localMem[1902]*7 + 6];
              ip = 4262;
      end

       4262 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[1913] == 0 ? 4292 : 4263;
      end

       4263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4263");
      end

       4264 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  4264");
      end

       4265 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4265");
      end

       4266 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  4266");
      end

       4267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4267");
      end

       4268 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4268");
      end

       4269 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4269");
      end

       4270 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4270");
      end

       4271 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4271");
      end

       4272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4272");
      end

       4273 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4273");
      end

       4274 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
         $display("Should not be executed  4274");
      end

       4275 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4275");
      end

       4276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4276");
      end

       4277 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4277");
      end

       4278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4278");
      end

       4279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4279");
      end

       4280 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4280");
      end

       4281 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4281");
      end

       4282 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4282");
      end

       4283 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4283");
      end

       4284 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  4284");
      end

       4285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4285");
      end

       4286 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4286");
      end

       4287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4287");
      end

       4288 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4288");
      end

       4289 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4289");
      end

       4290 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4290");
      end

       4291 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4291");
      end

       4292 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4293;
      end

       4293 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4294;
      end

       4294 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4295;
      end

       4295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1924] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4296;
      end

       4296 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4297;
      end

       4297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1926] = heapMem[localMem[1924]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4298;
      end

       4298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1927] = heapMem[localMem[1924]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4299;
      end

       4299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1928] = heapMem[localMem[1927]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4300;
      end

       4300 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[1926] <  localMem[1928] ? 4520 : 4301;
      end

       4301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4301");
      end

       4302 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  4302");
      end

       4303 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4303");
      end

       4304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4304");
      end

       4305 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4305");
      end

       4306 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4306");
      end

       4307 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4307");
      end

       4308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4308");
      end

       4309 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4309");
      end

       4310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4310");
      end

       4311 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4311");
      end

       4312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4312");
      end

       4313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4313");
      end

       4314 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4314");
      end

       4315 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4315");
      end

       4316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4316");
      end

       4317 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4317");
      end

       4318 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4318");
      end

       4319 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4319");
      end

       4320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4320");
      end

       4321 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4321");
      end

       4322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4322");
      end

       4323 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4323");
      end

       4324 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4324");
      end

       4325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4325");
      end

       4326 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4326");
      end

       4327 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4327");
      end

       4328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4328");
      end

       4329 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4329");
      end

       4330 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4330");
      end

       4331 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4331");
      end

       4332 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4332");
      end

       4333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4333");
      end

       4334 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4334");
      end

       4335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4335");
      end

       4336 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4336");
      end

       4337 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4337");
      end

       4338 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4338");
      end

       4339 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4339");
      end

       4340 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4340");
      end

       4341 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4341");
      end

       4342 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4342");
      end

       4343 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4343");
      end

       4344 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4344");
      end

       4345 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4345");
      end

       4346 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4346");
      end

       4347 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4347");
      end

       4348 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4348");
      end

       4349 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4349");
      end

       4350 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4350");
      end

       4351 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4351");
      end

       4352 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4352");
      end

       4353 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4353");
      end

       4354 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4354");
      end

       4355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4355");
      end

       4356 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4356");
      end

       4357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4357");
      end

       4358 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4358");
      end

       4359 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4359");
      end

       4360 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4360");
      end

       4361 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4361");
      end

       4362 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4362");
      end

       4363 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4363");
      end

       4364 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4364");
      end

       4365 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4365");
      end

       4366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4366");
      end

       4367 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4367");
      end

       4368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4368");
      end

       4369 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4369");
      end

       4370 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4370");
      end

       4371 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4371");
      end

       4372 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4372");
      end

       4373 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4373");
      end

       4374 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4374");
      end

       4375 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4375");
      end

       4376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4376");
      end

       4377 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4377");
      end

       4378 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4378");
      end

       4379 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4379");
      end

       4380 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  4380");
      end

       4381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4381");
      end

       4382 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  4382");
      end

       4383 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  4383");
      end

       4384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4384");
      end

       4385 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4385");
      end

       4386 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4386");
      end

       4387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4387");
      end

       4388 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4388");
      end

       4389 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4389");
      end

       4390 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4390");
      end

       4391 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4391");
      end

       4392 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4392");
      end

       4393 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4393");
      end

       4394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4394");
      end

       4395 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4395");
      end

       4396 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4396");
      end

       4397 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4397");
      end

       4398 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4398");
      end

       4399 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4399");
      end

       4400 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4400");
      end

       4401 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4401");
      end

       4402 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4402");
      end

       4403 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4403");
      end

       4404 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4404");
      end

       4405 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4405");
      end

       4406 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4406");
      end

       4407 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4407");
      end

       4408 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4408");
      end

       4409 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4409");
      end

       4410 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4410");
      end

       4411 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4411");
      end

       4412 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4412");
      end

       4413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4413");
      end

       4414 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4414");
      end

       4415 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4415");
      end

       4416 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4416");
      end

       4417 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4417");
      end

       4418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4418");
      end

       4419 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4419");
      end

       4420 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4420");
      end

       4421 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4421");
      end

       4422 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4422");
      end

       4423 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4423");
      end

       4424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4424");
      end

       4425 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4425");
      end

       4426 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4426");
      end

       4427 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4427");
      end

       4428 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4428");
      end

       4429 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4429");
      end

       4430 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4430");
      end

       4431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4431");
      end

       4432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4432");
      end

       4433 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4433");
      end

       4434 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4434");
      end

       4435 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4435");
      end

       4436 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4436");
      end

       4437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4437");
      end

       4438 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4438");
      end

       4439 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4439");
      end

       4440 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4440");
      end

       4441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4441");
      end

       4442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4442");
      end

       4443 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4443");
      end

       4444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4444");
      end

       4445 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4445");
      end

       4446 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4446");
      end

       4447 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4447");
      end

       4448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4448");
      end

       4449 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4449");
      end

       4450 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4450");
      end

       4451 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4451");
      end

       4452 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4452");
      end

       4453 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4453");
      end

       4454 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4454");
      end

       4455 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4455");
      end

       4456 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4456");
      end

       4457 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4457");
      end

       4458 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4458");
      end

       4459 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4459");
      end

       4460 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4460");
      end

       4461 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4461");
      end

       4462 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4462");
      end

       4463 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4463");
      end

       4464 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4464");
      end

       4465 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4465");
      end

       4466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4466");
      end

       4467 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4467");
      end

       4468 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4468");
      end

       4469 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4469");
      end

       4470 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4470");
      end

       4471 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4471");
      end

       4472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4472");
      end

       4473 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4473");
      end

       4474 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4474");
      end

       4475 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4475");
      end

       4476 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4476");
      end

       4477 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4477");
      end

       4478 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4478");
      end

       4479 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4479");
      end

       4480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4480");
      end

       4481 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4481");
      end

       4482 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4482");
      end

       4483 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4483");
      end

       4484 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4484");
      end

       4485 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4485");
      end

       4486 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4486");
      end

       4487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4487");
      end

       4488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4488");
      end

       4489 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4489");
      end

       4490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4490");
      end

       4491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4491");
      end

       4492 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4492");
      end

       4493 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4493");
      end

       4494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4494");
      end

       4495 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4495");
      end

       4496 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4496");
      end

       4497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4497");
      end

       4498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4498");
      end

       4499 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4499");
      end

       4500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4500");
      end

       4501 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4501");
      end

       4502 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4502");
      end

       4503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4503");
      end

       4504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4504");
      end

       4505 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4505");
      end

       4506 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4506");
      end

       4507 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4507");
      end

       4508 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4508");
      end

       4509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4509");
      end

       4510 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4510");
      end

       4511 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4511");
      end

       4512 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4512");
      end

       4513 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4513");
      end

       4514 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4514");
      end

       4515 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4515");
      end

       4516 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4516");
      end

       4517 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4517");
      end

       4518 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4518");
      end

       4519 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4519");
      end

       4520 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4521;
      end

       4521 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1925] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4522;
      end

       4522 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4523;
      end

       4523 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4524;
      end

       4524 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4525;
      end

       4525 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2032] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4526;
      end

       4526 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4527;
      end

       4527 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2032] >= 99 ? 5025 : 4528;
      end

       4528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2033] = heapMem[localMem[1924]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4529;
      end

       4529 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2034] = localMem[2033] - 1;
              updateArrayLength(2, 0, 0);
              ip = 4530;
      end

       4530 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2035] = heapMem[localMem[1924]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 4531;
      end

       4531 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2036] = heapMem[localMem[2035]*7 + localMem[2034]];
              updateArrayLength(2, 0, 0);
              ip = 4532;
      end

       4532 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 5 <= localMem[2036] ? 4773 : 4533;
      end

       4533 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2037] = !heapMem[localMem[1924]*7 + 6];
              ip = 4534;
      end

       4534 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2037] == 0 ? 4539 : 4535;
      end

       4535 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*7 + 0] = localMem[1924];
              updateArrayLength(1, localMem[1901], 0);
              ip = 4536;
      end

       4536 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[1901]*7 + 1] = 2;
              updateArrayLength(1, localMem[1901], 1);
              ip = 4537;
      end

       4537 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[1901]*7 + 2] = localMem[2033] - 1;
              updateArrayLength(1, localMem[1901], 2);
              ip = 4538;
      end

       4538 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5029;
      end

       4539 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4540;
      end

       4540 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2038] = heapMem[localMem[1924]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 4541;
      end

       4541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2039] = heapMem[localMem[2038]*7 + localMem[2033]];
              updateArrayLength(2, 0, 0);
              ip = 4542;
      end

       4542 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4543;
      end

       4543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2041] = heapMem[localMem[2039]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 4544;
      end

       4544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2042] = heapMem[localMem[2039]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 4545;
      end

       4545 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2043] = heapMem[localMem[2042]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 4546;
      end

       4546 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2041] <  localMem[2043] ? 4766 : 4547;
      end

       4547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4547");
      end

       4548 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  4548");
      end

       4549 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4549");
      end

       4550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4550");
      end

       4551 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4551");
      end

       4552 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4552");
      end

       4553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4553");
      end

       4554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4554");
      end

       4555 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4555");
      end

       4556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4556");
      end

       4557 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4557");
      end

       4558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4558");
      end

       4559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4559");
      end

       4560 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4560");
      end

       4561 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4561");
      end

       4562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4562");
      end

       4563 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4563");
      end

       4564 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4564");
      end

       4565 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4565");
      end

       4566 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4566");
      end

       4567 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4567");
      end

       4568 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4568");
      end

       4569 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4569");
      end

       4570 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4570");
      end

       4571 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4571");
      end

       4572 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4572");
      end

       4573 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4573");
      end

       4574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4574");
      end

       4575 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4575");
      end

       4576 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4576");
      end

       4577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4577");
      end

       4578 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4578");
      end

       4579 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4579");
      end

       4580 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4580");
      end

       4581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4581");
      end

       4582 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4582");
      end

       4583 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4583");
      end

       4584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4584");
      end

       4585 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4585");
      end

       4586 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4586");
      end

       4587 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4587");
      end

       4588 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4588");
      end

       4589 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4589");
      end

       4590 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4590");
      end

       4591 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4591");
      end

       4592 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4592");
      end

       4593 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4593");
      end

       4594 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4594");
      end

       4595 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4595");
      end

       4596 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4596");
      end

       4597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4597");
      end

       4598 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4598");
      end

       4599 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4599");
      end

       4600 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4600");
      end

       4601 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4601");
      end

       4602 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4602");
      end

       4603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4603");
      end

       4604 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4604");
      end

       4605 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4605");
      end

       4606 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4606");
      end

       4607 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4607");
      end

       4608 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4608");
      end

       4609 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4609");
      end

       4610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4610");
      end

       4611 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4611");
      end

       4612 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4612");
      end

       4613 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4613");
      end

       4614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4614");
      end

       4615 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4615");
      end

       4616 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4616");
      end

       4617 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4617");
      end

       4618 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4618");
      end

       4619 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4619");
      end

       4620 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4620");
      end

       4621 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4621");
      end

       4622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4622");
      end

       4623 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4623");
      end

       4624 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4624");
      end

       4625 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4625");
      end

       4626 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  4626");
      end

       4627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4627");
      end

       4628 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  4628");
      end

       4629 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  4629");
      end

       4630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4630");
      end

       4631 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4631");
      end

       4632 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4632");
      end

       4633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4633");
      end

       4634 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4634");
      end

       4635 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4635");
      end

       4636 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4636");
      end

       4637 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4637");
      end

       4638 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4638");
      end

       4639 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4639");
      end

       4640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4640");
      end

       4641 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4641");
      end

       4642 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4642");
      end

       4643 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4643");
      end

       4644 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4644");
      end

       4645 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4645");
      end

       4646 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4646");
      end

       4647 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4647");
      end

       4648 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4648");
      end

       4649 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4649");
      end

       4650 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4650");
      end

       4651 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4651");
      end

       4652 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4652");
      end

       4653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4653");
      end

       4654 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4654");
      end

       4655 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4655");
      end

       4656 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4656");
      end

       4657 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4657");
      end

       4658 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4658");
      end

       4659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4659");
      end

       4660 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4660");
      end

       4661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4661");
      end

       4662 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4662");
      end

       4663 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4663");
      end

       4664 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4664");
      end

       4665 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4665");
      end

       4666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4666");
      end

       4667 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4667");
      end

       4668 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4668");
      end

       4669 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4669");
      end

       4670 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4670");
      end

       4671 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4671");
      end

       4672 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4672");
      end

       4673 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4673");
      end

       4674 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4674");
      end

       4675 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4675");
      end

       4676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4676");
      end

       4677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4677");
      end

       4678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4678");
      end

       4679 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4679");
      end

       4680 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4680");
      end

       4681 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4681");
      end

       4682 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4682");
      end

       4683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4683");
      end

       4684 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4684");
      end

       4685 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4685");
      end

       4686 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4686");
      end

       4687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4687");
      end

       4688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4688");
      end

       4689 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4689");
      end

       4690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4690");
      end

       4691 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4691");
      end

       4692 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4692");
      end

       4693 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4693");
      end

       4694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4694");
      end

       4695 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4695");
      end

       4696 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4696");
      end

       4697 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4697");
      end

       4698 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4698");
      end

       4699 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4699");
      end

       4700 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4700");
      end

       4701 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4701");
      end

       4702 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4702");
      end

       4703 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4703");
      end

       4704 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4704");
      end

       4705 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4705");
      end

       4706 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4706");
      end

       4707 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4707");
      end

       4708 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4708");
      end

       4709 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4709");
      end

       4710 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4710");
      end

       4711 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4711");
      end

       4712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4712");
      end

       4713 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4713");
      end

       4714 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4714");
      end

       4715 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4715");
      end

       4716 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4716");
      end

       4717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4717");
      end

       4718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4718");
      end

       4719 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4719");
      end

       4720 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4720");
      end

       4721 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4721");
      end

       4722 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4722");
      end

       4723 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4723");
      end

       4724 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4724");
      end

       4725 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4725");
      end

       4726 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4726");
      end

       4727 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4727");
      end

       4728 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4728");
      end

       4729 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4729");
      end

       4730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4730");
      end

       4731 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4731");
      end

       4732 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4732");
      end

       4733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4733");
      end

       4734 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4734");
      end

       4735 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4735");
      end

       4736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4736");
      end

       4737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4737");
      end

       4738 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4738");
      end

       4739 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4739");
      end

       4740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4740");
      end

       4741 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4741");
      end

       4742 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4742");
      end

       4743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4743");
      end

       4744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4744");
      end

       4745 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4745");
      end

       4746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4746");
      end

       4747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4747");
      end

       4748 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4748");
      end

       4749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4749");
      end

       4750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4750");
      end

       4751 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4751");
      end

       4752 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4752");
      end

       4753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4753");
      end

       4754 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4754");
      end

       4755 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4755");
      end

       4756 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4756");
      end

       4757 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4757");
      end

       4758 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4758");
      end

       4759 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4759");
      end

       4760 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4760");
      end

       4761 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4761");
      end

       4762 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4762");
      end

       4763 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4763");
      end

       4764 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4764");
      end

       4765 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4765");
      end

       4766 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4767;
      end

       4767 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2040] = 0;
              updateArrayLength(2, 0, 0);
              ip = 4768;
      end

       4768 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4769;
      end

       4769 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2040] != 0 ? 4771 : 4770;
      end

       4770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[1924] = localMem[2039];
              updateArrayLength(2, 0, 0);
              ip = 4771;
      end

       4771 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 4772;
      end

       4772 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5022;
      end

       4773 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4773");
      end

       4774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4774");
      end

       4775 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  4775");
      end

       4776 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4776");
      end

       4777 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4777");
      end

       4778 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4778");
      end

       4779 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  4779");
      end

       4780 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4780");
      end

       4781 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4781");
      end

       4782 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  4782");
      end

       4783 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4783");
      end

       4784 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4784");
      end

       4785 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4785");
      end

       4786 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4786");
      end

       4787 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4787");
      end

       4788 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4788");
      end

       4789 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4789");
      end

       4790 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4790");
      end

       4791 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4791");
      end

       4792 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4792");
      end

       4793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4793");
      end

       4794 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4794");
      end

       4795 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4795");
      end

       4796 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  4796");
      end

       4797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4797");
      end

       4798 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  4798");
      end

       4799 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4799");
      end

       4800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4800");
      end

       4801 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  4801");
      end

       4802 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4802");
      end

       4803 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4803");
      end

       4804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4804");
      end

       4805 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4805");
      end

       4806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4806");
      end

       4807 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4807");
      end

       4808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4808");
      end

       4809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4809");
      end

       4810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4810");
      end

       4811 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4811");
      end

       4812 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4812");
      end

       4813 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4813");
      end

       4814 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4814");
      end

       4815 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4815");
      end

       4816 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4816");
      end

       4817 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4817");
      end

       4818 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4818");
      end

       4819 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4819");
      end

       4820 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4820");
      end

       4821 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4821");
      end

       4822 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4822");
      end

       4823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4823");
      end

       4824 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4824");
      end

       4825 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4825");
      end

       4826 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4826");
      end

       4827 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4827");
      end

       4828 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4828");
      end

       4829 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4829");
      end

       4830 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4830");
      end

       4831 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4831");
      end

       4832 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4832");
      end

       4833 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4833");
      end

       4834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4834");
      end

       4835 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4835");
      end

       4836 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4836");
      end

       4837 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4837");
      end

       4838 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4838");
      end

       4839 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4839");
      end

       4840 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4840");
      end

       4841 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4841");
      end

       4842 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4842");
      end

       4843 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4843");
      end

       4844 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4844");
      end

       4845 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4845");
      end

       4846 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4846");
      end

       4847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4847");
      end

       4848 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4848");
      end

       4849 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4849");
      end

       4850 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4850");
      end

       4851 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4851");
      end

       4852 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4852");
      end

       4853 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4853");
      end

       4854 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4854");
      end

       4855 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4855");
      end

       4856 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4856");
      end

       4857 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4857");
      end

       4858 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4858");
      end

       4859 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4859");
      end

       4860 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4860");
      end

       4861 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4861");
      end

       4862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4862");
      end

       4863 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4863");
      end

       4864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4864");
      end

       4865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4865");
      end

       4866 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4866");
      end

       4867 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4867");
      end

       4868 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4868");
      end

       4869 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4869");
      end

       4870 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4870");
      end

       4871 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4871");
      end

       4872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4872");
      end

       4873 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4873");
      end

       4874 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4874");
      end

       4875 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4875");
      end

       4876 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  4876");
      end

       4877 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4877");
      end

       4878 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  4878");
      end

       4879 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  4879");
      end

       4880 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4880");
      end

       4881 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4881");
      end

       4882 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4882");
      end

       4883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4883");
      end

       4884 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4884");
      end

       4885 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4885");
      end

       4886 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4886");
      end

       4887 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  4887");
      end

       4888 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4888");
      end

       4889 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4889");
      end

       4890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4890");
      end

       4891 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4891");
      end

       4892 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4892");
      end

       4893 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4893");
      end

       4894 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  4894");
      end

       4895 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4895");
      end

       4896 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4896");
      end

       4897 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4897");
      end

       4898 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4898");
      end

       4899 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4899");
      end

       4900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4900");
      end

       4901 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4901");
      end

       4902 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4902");
      end

       4903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4903");
      end

       4904 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4904");
      end

       4905 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4905");
      end

       4906 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4906");
      end

       4907 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4907");
      end

       4908 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4908");
      end

       4909 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4909");
      end

       4910 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4910");
      end

       4911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4911");
      end

       4912 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4912");
      end

       4913 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4913");
      end

       4914 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4914");
      end

       4915 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4915");
      end

       4916 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4916");
      end

       4917 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4917");
      end

       4918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4918");
      end

       4919 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4919");
      end

       4920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4920");
      end

       4921 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  4921");
      end

       4922 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  4922");
      end

       4923 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4923");
      end

       4924 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4924");
      end

       4925 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4925");
      end

       4926 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4926");
      end

       4927 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4927");
      end

       4928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4928");
      end

       4929 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4929");
      end

       4930 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4930");
      end

       4931 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4931");
      end

       4932 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4932");
      end

       4933 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4933");
      end

       4934 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4934");
      end

       4935 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4935");
      end

       4936 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4936");
      end

       4937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4937");
      end

       4938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4938");
      end

       4939 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4939");
      end

       4940 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4940");
      end

       4941 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4941");
      end

       4942 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4942");
      end

       4943 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4943");
      end

       4944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4944");
      end

       4945 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4945");
      end

       4946 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4946");
      end

       4947 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4947");
      end

       4948 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4948");
      end

       4949 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4949");
      end

       4950 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4950");
      end

       4951 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4951");
      end

       4952 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4952");
      end

       4953 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4953");
      end

       4954 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4954");
      end

       4955 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4955");
      end

       4956 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4956");
      end

       4957 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4957");
      end

       4958 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4958");
      end

       4959 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4959");
      end

       4960 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4960");
      end

       4961 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4961");
      end

       4962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4962");
      end

       4963 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4963");
      end

       4964 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4964");
      end

       4965 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4965");
      end

       4966 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  4966");
      end

       4967 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4967");
      end

       4968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4968");
      end

       4969 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4969");
      end

       4970 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  4970");
      end

       4971 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4971");
      end

       4972 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4972");
      end

       4973 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  4973");
      end

       4974 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4974");
      end

       4975 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  4975");
      end

       4976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4976");
      end

       4977 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4977");
      end

       4978 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4978");
      end

       4979 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4979");
      end

       4980 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4980");
      end

       4981 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4981");
      end

       4982 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4982");
      end

       4983 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4983");
      end

       4984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4984");
      end

       4985 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4985");
      end

       4986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4986");
      end

       4987 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4987");
      end

       4988 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  4988");
      end

       4989 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  4989");
      end

       4990 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4990");
      end

       4991 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4991");
      end

       4992 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4992");
      end

       4993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4993");
      end

       4994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4994");
      end

       4995 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4995");
      end

       4996 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4996");
      end

       4997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4997");
      end

       4998 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4998");
      end

       4999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  4999");
      end

       5000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5000");
      end

       5001 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5001");
      end

       5002 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5002");
      end

       5003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5003");
      end

       5004 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5004");
      end

       5005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5005");
      end

       5006 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5006");
      end

       5007 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5007");
      end

       5008 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5008");
      end

       5009 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5009");
      end

       5010 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5010");
      end

       5011 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5011");
      end

       5012 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5012");
      end

       5013 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5013");
      end

       5014 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5014");
      end

       5015 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5015");
      end

       5016 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5016");
      end

       5017 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5017");
      end

       5018 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5018");
      end

       5019 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5019");
      end

       5020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5020");
      end

       5021 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5021");
      end

       5022 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5023;
      end

       5023 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2032] = localMem[2032] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5024;
      end

       5024 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 4526;
      end

       5025 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5025");
      end

       5026 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
         $display("Should not be executed  5026");
      end

       5027 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5027");
      end

       5028 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5028");
      end

       5029 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5030;
      end

       5030 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2260] = heapMem[localMem[1901]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5031;
      end

       5031 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2261] = heapMem[localMem[1901]*7 + 1];
              updateArrayLength(2, 0, 0);
              ip = 5032;
      end

       5032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2262] = heapMem[localMem[1901]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5033;
      end

       5033 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2261] != 1 ? 5037 : 5034;
      end

       5034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5034");
      end

       5035 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5035");
      end

       5036 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5036");
      end

       5037 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5038;
      end

       5038 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2261] != 2 ? 5046 : 5039;
      end

       5039 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2264] = localMem[2262] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5040;
      end

       5040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2265] = heapMem[localMem[2260]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5041;
      end

       5041 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2265] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2264], localMem[2265], arraySizes[localMem[2265]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2264] && i <= arraySizes[localMem[2265]]) begin
                  heapMem[NArea * localMem[2265] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2265] + localMem[2264]] = 5;                                    // Insert new value
              arraySizes[localMem[2265]] = arraySizes[localMem[2265]] + 1;                              // Increase array size
              ip = 5042;
      end

       5042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2266] = heapMem[localMem[2260]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5043;
      end

       5043 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2266] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2264], localMem[2266], arraySizes[localMem[2266]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2264] && i <= arraySizes[localMem[2266]]) begin
                  heapMem[NArea * localMem[2266] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2266] + localMem[2264]] = 55;                                    // Insert new value
              arraySizes[localMem[2266]] = arraySizes[localMem[2266]] + 1;                              // Increase array size
              ip = 5044;
      end

       5044 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2260]*7 + 0] = heapMem[localMem[2260]*7 + 0] + 1;
              updateArrayLength(1, localMem[2260], 0);
              ip = 5045;
      end

       5045 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5052;
      end

       5046 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5046");
      end

       5047 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5047");
      end

       5048 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5048");
      end

       5049 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5049");
      end

       5050 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5050");
      end

       5051 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5051");
      end

       5052 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5053;
      end

       5053 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = heapMem[localMem[0]*7 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 5054;
      end

       5054 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5055;
      end

       5055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2270] = heapMem[localMem[2260]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5056;
      end

       5056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2271] = heapMem[localMem[2260]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5057;
      end

       5057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2272] = heapMem[localMem[2271]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5058;
      end

       5058 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2270] <  localMem[2272] ? 5278 : 5059;
      end

       5059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2273] = localMem[2272];
              updateArrayLength(2, 0, 0);
              ip = 5060;
      end

       5060 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
              localMem[2273] = localMem[2273] >> 1;
              ip = 5061;
      end

       5061 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2274] = localMem[2273] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5062;
      end

       5062 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2275] = heapMem[localMem[2260]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5063;
      end

       5063 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2275] == 0 ? 5160 : 5064;
      end

       5064 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2276] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2276] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2276]] = 0;
              ip = 5065;
      end

       5065 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 0] = localMem[2273];
              updateArrayLength(1, localMem[2276], 0);
              ip = 5066;
      end

       5066 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 2] = 0;
              updateArrayLength(1, localMem[2276], 2);
              ip = 5067;
      end

       5067 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2277] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2277] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2277]] = 0;
              ip = 5068;
      end

       5068 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 4] = localMem[2277];
              updateArrayLength(1, localMem[2276], 4);
              ip = 5069;
      end

       5069 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2278] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2278] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2278]] = 0;
              ip = 5070;
      end

       5070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 5] = localMem[2278];
              updateArrayLength(1, localMem[2276], 5);
              ip = 5071;
      end

       5071 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 6] = 0;
              updateArrayLength(1, localMem[2276], 6);
              ip = 5072;
      end

       5072 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 3] = localMem[2271];
              updateArrayLength(1, localMem[2276], 3);
              ip = 5073;
      end

       5073 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2271]*7 + 1] = heapMem[localMem[2271]*7 + 1] + 1;
              updateArrayLength(1, localMem[2271], 1);
              ip = 5074;
      end

       5074 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 1] = heapMem[localMem[2271]*7 + 1];
              updateArrayLength(1, localMem[2276], 1);
              ip = 5075;
      end

       5075 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2279] = !heapMem[localMem[2260]*7 + 6];
              ip = 5076;
      end

       5076 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2279] != 0 ? 5105 : 5077;
      end

       5077 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5077");
      end

       5078 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5078");
      end

       5079 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5079");
      end

       5080 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5080");
      end

       5081 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5081");
      end

       5082 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5082");
      end

       5083 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5083");
      end

       5084 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5084");
      end

       5085 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5085");
      end

       5086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5086");
      end

       5087 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5087");
      end

       5088 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5088");
      end

       5089 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5089");
      end

       5090 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5090");
      end

       5091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5091");
      end

       5092 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5092");
      end

       5093 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5093");
      end

       5094 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5094");
      end

       5095 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5095");
      end

       5096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5096");
      end

       5097 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5097");
      end

       5098 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5098");
      end

       5099 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5099");
      end

       5100 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5100");
      end

       5101 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5101");
      end

       5102 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5102");
      end

       5103 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5103");
      end

       5104 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5104");
      end

       5105 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5106;
      end

       5106 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2294] = heapMem[localMem[2260]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5107;
      end

       5107 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2295] = heapMem[localMem[2276]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5108;
      end

       5108 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2295] + 0 + i] = heapMem[NArea * localMem[2294] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2295], 0 + i);
                end
              end
              ip = 5109;
      end

       5109 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2296] = heapMem[localMem[2260]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5110;
      end

       5110 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2297] = heapMem[localMem[2276]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5111;
      end

       5111 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
              for(i = 0; i < NArea; i = i + 1) begin                            // Copy from source to target
                if (i < localMem[2273]) begin
                  heapMem[NArea * localMem[2297] + 0 + i] = heapMem[NArea * localMem[2296] + localMem[2274] + i];
                  updateArrayLength(1, localMem[2297], 0 + i);
                end
              end
              ip = 5112;
      end

       5112 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5113;
      end

       5113 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2260]*7 + 0] = localMem[2273];
              updateArrayLength(1, localMem[2260], 0);
              ip = 5114;
      end

       5114 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2276]*7 + 2] = localMem[2275];
              updateArrayLength(1, localMem[2276], 2);
              ip = 5115;
      end

       5115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2298] = heapMem[localMem[2275]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5116;
      end

       5116 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2299] = heapMem[localMem[2275]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5117;
      end

       5117 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2300] = heapMem[localMem[2299]*7 + localMem[2298]];
              updateArrayLength(2, 0, 0);
              ip = 5118;
      end

       5118 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2300] != localMem[2260] ? 5137 : 5119;
      end

       5119 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2301] = heapMem[localMem[2260]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5120;
      end

       5120 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2302] = heapMem[localMem[2301]*7 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5121;
      end

       5121 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2303] = heapMem[localMem[2275]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5122;
      end

       5122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2303]*7 + localMem[2298]] = localMem[2302];
              updateArrayLength(1, localMem[2303], localMem[2298]);
              ip = 5123;
      end

       5123 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2304] = heapMem[localMem[2260]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5124;
      end

       5124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2305] = heapMem[localMem[2304]*7 + localMem[2273]];
              updateArrayLength(2, 0, 0);
              ip = 5125;
      end

       5125 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2306] = heapMem[localMem[2275]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5126;
      end

       5126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2306]*7 + localMem[2298]] = localMem[2305];
              updateArrayLength(1, localMem[2306], localMem[2298]);
              ip = 5127;
      end

       5127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2307] = heapMem[localMem[2260]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5128;
      end

       5128 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2307]] = localMem[2273];
              ip = 5129;
      end

       5129 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2308] = heapMem[localMem[2260]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 5130;
      end

       5130 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
              arraySizes[localMem[2308]] = localMem[2273];
              ip = 5131;
      end

       5131 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2309] = localMem[2298] + 1;
              updateArrayLength(2, 0, 0);
              ip = 5132;
      end

       5132 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2275]*7 + 0] = localMem[2309];
              updateArrayLength(1, localMem[2275], 0);
              ip = 5133;
      end

       5133 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2310] = heapMem[localMem[2275]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5134;
      end

       5134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2310]*7 + localMem[2309]] = localMem[2276];
              updateArrayLength(1, localMem[2310], localMem[2309]);
              ip = 5135;
      end

       5135 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5275;
      end

       5136 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5136");
      end

       5137 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5137");
      end

       5138 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  5138");
      end

       5139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5139");
      end

       5140 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  5140");
      end

       5141 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  5141");
      end

       5142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5142");
      end

       5143 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5143");
      end

       5144 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5144");
      end

       5145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5145");
      end

       5146 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5146");
      end

       5147 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5147");
      end

       5148 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5148");
      end

       5149 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5149");
      end

       5150 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5150");
      end

       5151 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5151");
      end

       5152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5152");
      end

       5153 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5153");
      end

       5154 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5154");
      end

       5155 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5155");
      end

       5156 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5156");
      end

       5157 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5157");
      end

       5158 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5158");
      end

       5159 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5159");
      end

       5160 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5160");
      end

       5161 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5161");
      end

       5162 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5162");
      end

       5163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5163");
      end

       5164 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5164");
      end

       5165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5165");
      end

       5166 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5166");
      end

       5167 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5167");
      end

       5168 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5168");
      end

       5169 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5169");
      end

       5170 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5170");
      end

       5171 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5171");
      end

       5172 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5172");
      end

       5173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5173");
      end

       5174 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5174");
      end

       5175 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5175");
      end

       5176 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5176");
      end

       5177 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5177");
      end

       5178 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5178");
      end

       5179 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5179");
      end

       5180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5180");
      end

       5181 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5181");
      end

       5182 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5182");
      end

       5183 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5183");
      end

       5184 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5184");
      end

       5185 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5185");
      end

       5186 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5186");
      end

       5187 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5187");
      end

       5188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5188");
      end

       5189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5189");
      end

       5190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5190");
      end

       5191 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5191");
      end

       5192 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5192");
      end

       5193 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5193");
      end

       5194 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5194");
      end

       5195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5195");
      end

       5196 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5196");
      end

       5197 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5197");
      end

       5198 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5198");
      end

       5199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5199");
      end

       5200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5200");
      end

       5201 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5201");
      end

       5202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5202");
      end

       5203 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5203");
      end

       5204 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5204");
      end

       5205 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5205");
      end

       5206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5206");
      end

       5207 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5207");
      end

       5208 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5208");
      end

       5209 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5209");
      end

       5210 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5210");
      end

       5211 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5211");
      end

       5212 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5212");
      end

       5213 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5213");
      end

       5214 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5214");
      end

       5215 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5215");
      end

       5216 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5216");
      end

       5217 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5217");
      end

       5218 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5218");
      end

       5219 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5219");
      end

       5220 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5220");
      end

       5221 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5221");
      end

       5222 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5222");
      end

       5223 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5223");
      end

       5224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5224");
      end

       5225 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5225");
      end

       5226 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5226");
      end

       5227 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5227");
      end

       5228 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5228");
      end

       5229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5229");
      end

       5230 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5230");
      end

       5231 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5231");
      end

       5232 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5232");
      end

       5233 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5233");
      end

       5234 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5234");
      end

       5235 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5235");
      end

       5236 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5236");
      end

       5237 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5237");
      end

       5238 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5238");
      end

       5239 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5239");
      end

       5240 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5240");
      end

       5241 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5241");
      end

       5242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5242");
      end

       5243 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5243");
      end

       5244 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5244");
      end

       5245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5245");
      end

       5246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5246");
      end

       5247 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5247");
      end

       5248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5248");
      end

       5249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5249");
      end

       5250 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5250");
      end

       5251 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5251");
      end

       5252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5252");
      end

       5253 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5253");
      end

       5254 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5254");
      end

       5255 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5255");
      end

       5256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5256");
      end

       5257 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5257");
      end

       5258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5258");
      end

       5259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5259");
      end

       5260 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5260");
      end

       5261 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5261");
      end

       5262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5262");
      end

       5263 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5263");
      end

       5264 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5264");
      end

       5265 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5265");
      end

       5266 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5266");
      end

       5267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5267");
      end

       5268 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5268");
      end

       5269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5269");
      end

       5270 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5270");
      end

       5271 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5271");
      end

       5272 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5272");
      end

       5273 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5273");
      end

       5274 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5274");
      end

       5275 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5276;
      end

       5276 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2269] = 1;
              updateArrayLength(2, 0, 0);
              ip = 5277;
      end

       5277 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5280;
      end

       5278 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5278");
      end

       5279 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5279");
      end

       5280 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5281;
      end

       5281 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5282;
      end

       5282 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5283;
      end

       5283 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5284;
      end

       5284 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[1901]] = 0;
              freedArrays[freedArraysTop] = localMem[1901];
              freedArraysTop = freedArraysTop + 1;
              ip = 5285;
      end

       5285 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
              if (freedArraysTop > 0) begin
                freedArraysTop = freedArraysTop - 1;
                localMem[2376] = freedArrays[freedArraysTop];
              end
              else begin
                localMem[2376] = allocs;
                allocs = allocs + 1;

              end
              arraySizes[localMem[2376]] = 0;
              ip = 5286;
      end

       5286 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5287;
      end

       5287 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2377] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5288;
      end

       5288 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2377] != 0 ? 5311 : 5289;
      end

       5289 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5289");
      end

       5290 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5290");
      end

       5291 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5291");
      end

       5292 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5292");
      end

       5293 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5293");
      end

       5294 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5294");
      end

       5295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5295");
      end

       5296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5296");
      end

       5297 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5297");
      end

       5298 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5298");
      end

       5299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5299");
      end

       5300 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5300");
      end

       5301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5301");
      end

       5302 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5302");
      end

       5303 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5303");
      end

       5304 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5304");
      end

       5305 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5305");
      end

       5306 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5306");
      end

       5307 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5307");
      end

       5308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5308");
      end

       5309 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5309");
      end

       5310 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5310");
      end

       5311 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5312;
      end

       5312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2385] = heapMem[localMem[2377]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5313;
      end

       5313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2386] = heapMem[localMem[0]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5314;
      end

       5314 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2385] >= localMem[2386] ? 5350 : 5315;
      end

       5315 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2387] = heapMem[localMem[2377]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5316;
      end

       5316 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2387] != 0 ? 5349 : 5317;
      end

       5317 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2388] = !heapMem[localMem[2377]*7 + 6];
              ip = 5318;
      end

       5318 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2388] == 0 ? 5348 : 5319;
      end

       5319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5319");
      end

       5320 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  5320");
      end

       5321 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  5321");
      end

       5322 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  5322");
      end

       5323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5323");
      end

       5324 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5324");
      end

       5325 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5325");
      end

       5326 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5326");
      end

       5327 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5327");
      end

       5328 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5328");
      end

       5329 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5329");
      end

       5330 :
      begin                                                                     // arrayCountGreater
if (0) begin
  $display("AAAA %4d %4d arrayCountGreater", steps, ip);
end
         $display("Should not be executed  5330");
      end

       5331 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5331");
      end

       5332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5332");
      end

       5333 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5333");
      end

       5334 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5334");
      end

       5335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5335");
      end

       5336 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5336");
      end

       5337 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5337");
      end

       5338 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5338");
      end

       5339 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5339");
      end

       5340 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  5340");
      end

       5341 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5341");
      end

       5342 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5342");
      end

       5343 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5343");
      end

       5344 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5344");
      end

       5345 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5345");
      end

       5346 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5346");
      end

       5347 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5347");
      end

       5348 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5349;
      end

       5349 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5350;
      end

       5350 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5351;
      end

       5351 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2399] = heapMem[localMem[0]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5352;
      end

       5352 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5353;
      end

       5353 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2401] = heapMem[localMem[2399]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5354;
      end

       5354 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2402] = heapMem[localMem[2399]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5355;
      end

       5355 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2403] = heapMem[localMem[2402]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5356;
      end

       5356 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2401] <  localMem[2403] ? 5576 : 5357;
      end

       5357 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5357");
      end

       5358 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  5358");
      end

       5359 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5359");
      end

       5360 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5360");
      end

       5361 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  5361");
      end

       5362 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5362");
      end

       5363 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5363");
      end

       5364 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5364");
      end

       5365 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5365");
      end

       5366 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5366");
      end

       5367 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5367");
      end

       5368 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5368");
      end

       5369 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5369");
      end

       5370 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5370");
      end

       5371 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5371");
      end

       5372 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5372");
      end

       5373 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5373");
      end

       5374 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5374");
      end

       5375 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5375");
      end

       5376 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5376");
      end

       5377 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5377");
      end

       5378 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5378");
      end

       5379 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5379");
      end

       5380 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5380");
      end

       5381 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5381");
      end

       5382 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5382");
      end

       5383 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5383");
      end

       5384 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5384");
      end

       5385 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5385");
      end

       5386 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5386");
      end

       5387 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5387");
      end

       5388 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5388");
      end

       5389 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5389");
      end

       5390 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5390");
      end

       5391 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5391");
      end

       5392 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5392");
      end

       5393 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5393");
      end

       5394 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5394");
      end

       5395 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5395");
      end

       5396 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5396");
      end

       5397 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5397");
      end

       5398 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5398");
      end

       5399 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5399");
      end

       5400 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5400");
      end

       5401 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5401");
      end

       5402 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5402");
      end

       5403 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5403");
      end

       5404 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5404");
      end

       5405 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5405");
      end

       5406 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5406");
      end

       5407 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5407");
      end

       5408 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5408");
      end

       5409 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5409");
      end

       5410 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5410");
      end

       5411 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5411");
      end

       5412 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5412");
      end

       5413 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5413");
      end

       5414 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5414");
      end

       5415 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5415");
      end

       5416 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5416");
      end

       5417 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5417");
      end

       5418 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5418");
      end

       5419 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5419");
      end

       5420 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5420");
      end

       5421 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5421");
      end

       5422 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5422");
      end

       5423 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5423");
      end

       5424 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5424");
      end

       5425 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5425");
      end

       5426 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5426");
      end

       5427 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5427");
      end

       5428 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5428");
      end

       5429 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5429");
      end

       5430 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5430");
      end

       5431 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5431");
      end

       5432 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5432");
      end

       5433 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5433");
      end

       5434 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5434");
      end

       5435 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5435");
      end

       5436 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  5436");
      end

       5437 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5437");
      end

       5438 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  5438");
      end

       5439 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  5439");
      end

       5440 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5440");
      end

       5441 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5441");
      end

       5442 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5442");
      end

       5443 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5443");
      end

       5444 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5444");
      end

       5445 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5445");
      end

       5446 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5446");
      end

       5447 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5447");
      end

       5448 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5448");
      end

       5449 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5449");
      end

       5450 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5450");
      end

       5451 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5451");
      end

       5452 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5452");
      end

       5453 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5453");
      end

       5454 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5454");
      end

       5455 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5455");
      end

       5456 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5456");
      end

       5457 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5457");
      end

       5458 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5458");
      end

       5459 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5459");
      end

       5460 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5460");
      end

       5461 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5461");
      end

       5462 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5462");
      end

       5463 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5463");
      end

       5464 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5464");
      end

       5465 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5465");
      end

       5466 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5466");
      end

       5467 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5467");
      end

       5468 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5468");
      end

       5469 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5469");
      end

       5470 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5470");
      end

       5471 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5471");
      end

       5472 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5472");
      end

       5473 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5473");
      end

       5474 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5474");
      end

       5475 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5475");
      end

       5476 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5476");
      end

       5477 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5477");
      end

       5478 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5478");
      end

       5479 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5479");
      end

       5480 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5480");
      end

       5481 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5481");
      end

       5482 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5482");
      end

       5483 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5483");
      end

       5484 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5484");
      end

       5485 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5485");
      end

       5486 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5486");
      end

       5487 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5487");
      end

       5488 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5488");
      end

       5489 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5489");
      end

       5490 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5490");
      end

       5491 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5491");
      end

       5492 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5492");
      end

       5493 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5493");
      end

       5494 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5494");
      end

       5495 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5495");
      end

       5496 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5496");
      end

       5497 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5497");
      end

       5498 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5498");
      end

       5499 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5499");
      end

       5500 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5500");
      end

       5501 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5501");
      end

       5502 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5502");
      end

       5503 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5503");
      end

       5504 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5504");
      end

       5505 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5505");
      end

       5506 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5506");
      end

       5507 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5507");
      end

       5508 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5508");
      end

       5509 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5509");
      end

       5510 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5510");
      end

       5511 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5511");
      end

       5512 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5512");
      end

       5513 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5513");
      end

       5514 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5514");
      end

       5515 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5515");
      end

       5516 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5516");
      end

       5517 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5517");
      end

       5518 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5518");
      end

       5519 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5519");
      end

       5520 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5520");
      end

       5521 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5521");
      end

       5522 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5522");
      end

       5523 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5523");
      end

       5524 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5524");
      end

       5525 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5525");
      end

       5526 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5526");
      end

       5527 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5527");
      end

       5528 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5528");
      end

       5529 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5529");
      end

       5530 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5530");
      end

       5531 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5531");
      end

       5532 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5532");
      end

       5533 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5533");
      end

       5534 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5534");
      end

       5535 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5535");
      end

       5536 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5536");
      end

       5537 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5537");
      end

       5538 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5538");
      end

       5539 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5539");
      end

       5540 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5540");
      end

       5541 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5541");
      end

       5542 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5542");
      end

       5543 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5543");
      end

       5544 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5544");
      end

       5545 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5545");
      end

       5546 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5546");
      end

       5547 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5547");
      end

       5548 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5548");
      end

       5549 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5549");
      end

       5550 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5550");
      end

       5551 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5551");
      end

       5552 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5552");
      end

       5553 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5553");
      end

       5554 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5554");
      end

       5555 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5555");
      end

       5556 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5556");
      end

       5557 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5557");
      end

       5558 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5558");
      end

       5559 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5559");
      end

       5560 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5560");
      end

       5561 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5561");
      end

       5562 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5562");
      end

       5563 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5563");
      end

       5564 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5564");
      end

       5565 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5565");
      end

       5566 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5566");
      end

       5567 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5567");
      end

       5568 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5568");
      end

       5569 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5569");
      end

       5570 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5570");
      end

       5571 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5571");
      end

       5572 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5572");
      end

       5573 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5573");
      end

       5574 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5574");
      end

       5575 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5575");
      end

       5576 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5577;
      end

       5577 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2400] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5578;
      end

       5578 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5579;
      end

       5579 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5580;
      end

       5580 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5581;
      end

       5581 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2507] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5582;
      end

       5582 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5583;
      end

       5583 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
              ip = localMem[2507] >= 99 ? 6081 : 5584;
      end

       5584 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2508] = heapMem[localMem[2399]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5585;
      end

       5585 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              localMem[2509] = localMem[2508] - 1;
              updateArrayLength(2, 0, 0);
              ip = 5586;
      end

       5586 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2510] = heapMem[localMem[2399]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 5587;
      end

       5587 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2511] = heapMem[localMem[2510]*7 + localMem[2509]];
              updateArrayLength(2, 0, 0);
              ip = 5588;
      end

       5588 :
      begin                                                                     // jLe
if (0) begin
  $display("AAAA %4d %4d jLe", steps, ip);
end
              ip = 6 <= localMem[2511] ? 5829 : 5589;
      end

       5589 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
              localMem[2512] = !heapMem[localMem[2399]*7 + 6];
              ip = 5590;
      end

       5590 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
              ip = localMem[2512] == 0 ? 5595 : 5591;
      end

       5591 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*7 + 0] = localMem[2399];
              updateArrayLength(1, localMem[2376], 0);
              ip = 5592;
      end

       5592 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              heapMem[localMem[2376]*7 + 1] = 2;
              updateArrayLength(1, localMem[2376], 1);
              ip = 5593;
      end

       5593 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
              heapMem[localMem[2376]*7 + 2] = localMem[2508] - 1;
              updateArrayLength(1, localMem[2376], 2);
              ip = 5594;
      end

       5594 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6085;
      end

       5595 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5596;
      end

       5596 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2513] = heapMem[localMem[2399]*7 + 6];
              updateArrayLength(2, 0, 0);
              ip = 5597;
      end

       5597 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2514] = heapMem[localMem[2513]*7 + localMem[2508]];
              updateArrayLength(2, 0, 0);
              ip = 5598;
      end

       5598 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5599;
      end

       5599 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2516] = heapMem[localMem[2514]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 5600;
      end

       5600 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2517] = heapMem[localMem[2514]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 5601;
      end

       5601 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2518] = heapMem[localMem[2517]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 5602;
      end

       5602 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2516] <  localMem[2518] ? 5822 : 5603;
      end

       5603 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5603");
      end

       5604 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  5604");
      end

       5605 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5605");
      end

       5606 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5606");
      end

       5607 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  5607");
      end

       5608 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5608");
      end

       5609 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5609");
      end

       5610 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5610");
      end

       5611 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5611");
      end

       5612 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5612");
      end

       5613 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5613");
      end

       5614 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5614");
      end

       5615 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5615");
      end

       5616 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5616");
      end

       5617 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5617");
      end

       5618 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5618");
      end

       5619 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5619");
      end

       5620 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5620");
      end

       5621 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5621");
      end

       5622 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5622");
      end

       5623 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5623");
      end

       5624 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5624");
      end

       5625 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5625");
      end

       5626 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5626");
      end

       5627 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5627");
      end

       5628 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5628");
      end

       5629 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5629");
      end

       5630 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5630");
      end

       5631 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5631");
      end

       5632 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5632");
      end

       5633 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5633");
      end

       5634 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5634");
      end

       5635 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5635");
      end

       5636 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5636");
      end

       5637 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5637");
      end

       5638 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5638");
      end

       5639 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5639");
      end

       5640 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5640");
      end

       5641 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5641");
      end

       5642 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5642");
      end

       5643 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5643");
      end

       5644 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5644");
      end

       5645 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5645");
      end

       5646 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5646");
      end

       5647 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5647");
      end

       5648 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5648");
      end

       5649 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5649");
      end

       5650 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5650");
      end

       5651 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5651");
      end

       5652 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5652");
      end

       5653 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5653");
      end

       5654 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5654");
      end

       5655 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5655");
      end

       5656 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5656");
      end

       5657 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5657");
      end

       5658 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5658");
      end

       5659 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5659");
      end

       5660 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5660");
      end

       5661 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5661");
      end

       5662 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5662");
      end

       5663 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5663");
      end

       5664 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5664");
      end

       5665 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5665");
      end

       5666 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5666");
      end

       5667 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5667");
      end

       5668 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5668");
      end

       5669 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5669");
      end

       5670 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5670");
      end

       5671 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5671");
      end

       5672 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5672");
      end

       5673 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5673");
      end

       5674 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5674");
      end

       5675 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5675");
      end

       5676 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5676");
      end

       5677 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5677");
      end

       5678 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5678");
      end

       5679 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5679");
      end

       5680 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5680");
      end

       5681 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5681");
      end

       5682 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  5682");
      end

       5683 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5683");
      end

       5684 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  5684");
      end

       5685 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  5685");
      end

       5686 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5686");
      end

       5687 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5687");
      end

       5688 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5688");
      end

       5689 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5689");
      end

       5690 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5690");
      end

       5691 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5691");
      end

       5692 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5692");
      end

       5693 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5693");
      end

       5694 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5694");
      end

       5695 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5695");
      end

       5696 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5696");
      end

       5697 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5697");
      end

       5698 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5698");
      end

       5699 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5699");
      end

       5700 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5700");
      end

       5701 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5701");
      end

       5702 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5702");
      end

       5703 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5703");
      end

       5704 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5704");
      end

       5705 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5705");
      end

       5706 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5706");
      end

       5707 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5707");
      end

       5708 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5708");
      end

       5709 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5709");
      end

       5710 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5710");
      end

       5711 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5711");
      end

       5712 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5712");
      end

       5713 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5713");
      end

       5714 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5714");
      end

       5715 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5715");
      end

       5716 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5716");
      end

       5717 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5717");
      end

       5718 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5718");
      end

       5719 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5719");
      end

       5720 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5720");
      end

       5721 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5721");
      end

       5722 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5722");
      end

       5723 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5723");
      end

       5724 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5724");
      end

       5725 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5725");
      end

       5726 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5726");
      end

       5727 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5727");
      end

       5728 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5728");
      end

       5729 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5729");
      end

       5730 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5730");
      end

       5731 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5731");
      end

       5732 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5732");
      end

       5733 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5733");
      end

       5734 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5734");
      end

       5735 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5735");
      end

       5736 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5736");
      end

       5737 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5737");
      end

       5738 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5738");
      end

       5739 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5739");
      end

       5740 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5740");
      end

       5741 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5741");
      end

       5742 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5742");
      end

       5743 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5743");
      end

       5744 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5744");
      end

       5745 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5745");
      end

       5746 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5746");
      end

       5747 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5747");
      end

       5748 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5748");
      end

       5749 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5749");
      end

       5750 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5750");
      end

       5751 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5751");
      end

       5752 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5752");
      end

       5753 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5753");
      end

       5754 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5754");
      end

       5755 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5755");
      end

       5756 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5756");
      end

       5757 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5757");
      end

       5758 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5758");
      end

       5759 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5759");
      end

       5760 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5760");
      end

       5761 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5761");
      end

       5762 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5762");
      end

       5763 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5763");
      end

       5764 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5764");
      end

       5765 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5765");
      end

       5766 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5766");
      end

       5767 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5767");
      end

       5768 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5768");
      end

       5769 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5769");
      end

       5770 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5770");
      end

       5771 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5771");
      end

       5772 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5772");
      end

       5773 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5773");
      end

       5774 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5774");
      end

       5775 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5775");
      end

       5776 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5776");
      end

       5777 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5777");
      end

       5778 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5778");
      end

       5779 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5779");
      end

       5780 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5780");
      end

       5781 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5781");
      end

       5782 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5782");
      end

       5783 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5783");
      end

       5784 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5784");
      end

       5785 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5785");
      end

       5786 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5786");
      end

       5787 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5787");
      end

       5788 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5788");
      end

       5789 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5789");
      end

       5790 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5790");
      end

       5791 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5791");
      end

       5792 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5792");
      end

       5793 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5793");
      end

       5794 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5794");
      end

       5795 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5795");
      end

       5796 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5796");
      end

       5797 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5797");
      end

       5798 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5798");
      end

       5799 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5799");
      end

       5800 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5800");
      end

       5801 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5801");
      end

       5802 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5802");
      end

       5803 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5803");
      end

       5804 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5804");
      end

       5805 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5805");
      end

       5806 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5806");
      end

       5807 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5807");
      end

       5808 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5808");
      end

       5809 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5809");
      end

       5810 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5810");
      end

       5811 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5811");
      end

       5812 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5812");
      end

       5813 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5813");
      end

       5814 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5814");
      end

       5815 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5815");
      end

       5816 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5816");
      end

       5817 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5817");
      end

       5818 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5818");
      end

       5819 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5819");
      end

       5820 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5820");
      end

       5821 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5821");
      end

       5822 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5823;
      end

       5823 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2515] = 0;
              updateArrayLength(2, 0, 0);
              ip = 5824;
      end

       5824 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5825;
      end

       5825 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2515] != 0 ? 5827 : 5826;
      end

       5826 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2399] = localMem[2514];
              updateArrayLength(2, 0, 0);
              ip = 5827;
      end

       5827 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 5828;
      end

       5828 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6078;
      end

       5829 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5829");
      end

       5830 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5830");
      end

       5831 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  5831");
      end

       5832 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  5832");
      end

       5833 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5833");
      end

       5834 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5834");
      end

       5835 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  5835");
      end

       5836 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5836");
      end

       5837 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5837");
      end

       5838 :
      begin                                                                     // arrayCountLess
if (0) begin
  $display("AAAA %4d %4d arrayCountLess", steps, ip);
end
         $display("Should not be executed  5838");
      end

       5839 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5839");
      end

       5840 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  5840");
      end

       5841 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5841");
      end

       5842 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5842");
      end

       5843 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5843");
      end

       5844 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5844");
      end

       5845 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5845");
      end

       5846 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5846");
      end

       5847 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5847");
      end

       5848 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5848");
      end

       5849 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5849");
      end

       5850 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5850");
      end

       5851 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5851");
      end

       5852 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
         $display("Should not be executed  5852");
      end

       5853 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5853");
      end

       5854 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  5854");
      end

       5855 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5855");
      end

       5856 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5856");
      end

       5857 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  5857");
      end

       5858 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5858");
      end

       5859 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5859");
      end

       5860 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5860");
      end

       5861 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5861");
      end

       5862 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5862");
      end

       5863 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5863");
      end

       5864 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5864");
      end

       5865 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5865");
      end

       5866 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5866");
      end

       5867 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5867");
      end

       5868 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5868");
      end

       5869 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5869");
      end

       5870 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5870");
      end

       5871 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5871");
      end

       5872 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5872");
      end

       5873 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5873");
      end

       5874 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5874");
      end

       5875 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5875");
      end

       5876 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5876");
      end

       5877 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5877");
      end

       5878 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5878");
      end

       5879 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5879");
      end

       5880 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5880");
      end

       5881 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5881");
      end

       5882 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5882");
      end

       5883 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5883");
      end

       5884 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5884");
      end

       5885 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5885");
      end

       5886 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5886");
      end

       5887 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5887");
      end

       5888 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5888");
      end

       5889 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  5889");
      end

       5890 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5890");
      end

       5891 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5891");
      end

       5892 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5892");
      end

       5893 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5893");
      end

       5894 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5894");
      end

       5895 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5895");
      end

       5896 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5896");
      end

       5897 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5897");
      end

       5898 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5898");
      end

       5899 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5899");
      end

       5900 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5900");
      end

       5901 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5901");
      end

       5902 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5902");
      end

       5903 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5903");
      end

       5904 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5904");
      end

       5905 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5905");
      end

       5906 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5906");
      end

       5907 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5907");
      end

       5908 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5908");
      end

       5909 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5909");
      end

       5910 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5910");
      end

       5911 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5911");
      end

       5912 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5912");
      end

       5913 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5913");
      end

       5914 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5914");
      end

       5915 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5915");
      end

       5916 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5916");
      end

       5917 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5917");
      end

       5918 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5918");
      end

       5919 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5919");
      end

       5920 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5920");
      end

       5921 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5921");
      end

       5922 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5922");
      end

       5923 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5923");
      end

       5924 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5924");
      end

       5925 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5925");
      end

       5926 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5926");
      end

       5927 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5927");
      end

       5928 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5928");
      end

       5929 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5929");
      end

       5930 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5930");
      end

       5931 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5931");
      end

       5932 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  5932");
      end

       5933 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5933");
      end

       5934 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  5934");
      end

       5935 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  5935");
      end

       5936 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5936");
      end

       5937 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5937");
      end

       5938 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5938");
      end

       5939 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5939");
      end

       5940 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5940");
      end

       5941 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5941");
      end

       5942 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5942");
      end

       5943 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  5943");
      end

       5944 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5944");
      end

       5945 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5945");
      end

       5946 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5946");
      end

       5947 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5947");
      end

       5948 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5948");
      end

       5949 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5949");
      end

       5950 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  5950");
      end

       5951 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5951");
      end

       5952 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  5952");
      end

       5953 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5953");
      end

       5954 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  5954");
      end

       5955 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5955");
      end

       5956 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5956");
      end

       5957 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5957");
      end

       5958 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5958");
      end

       5959 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5959");
      end

       5960 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5960");
      end

       5961 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5961");
      end

       5962 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5962");
      end

       5963 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5963");
      end

       5964 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5964");
      end

       5965 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5965");
      end

       5966 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5966");
      end

       5967 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5967");
      end

       5968 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5968");
      end

       5969 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5969");
      end

       5970 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5970");
      end

       5971 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5971");
      end

       5972 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5972");
      end

       5973 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5973");
      end

       5974 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5974");
      end

       5975 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5975");
      end

       5976 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5976");
      end

       5977 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  5977");
      end

       5978 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  5978");
      end

       5979 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5979");
      end

       5980 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5980");
      end

       5981 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  5981");
      end

       5982 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5982");
      end

       5983 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5983");
      end

       5984 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5984");
      end

       5985 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5985");
      end

       5986 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5986");
      end

       5987 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5987");
      end

       5988 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5988");
      end

       5989 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5989");
      end

       5990 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5990");
      end

       5991 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  5991");
      end

       5992 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5992");
      end

       5993 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5993");
      end

       5994 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5994");
      end

       5995 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5995");
      end

       5996 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5996");
      end

       5997 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5997");
      end

       5998 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  5998");
      end

       5999 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  5999");
      end

       6000 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6000");
      end

       6001 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6001");
      end

       6002 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6002");
      end

       6003 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6003");
      end

       6004 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6004");
      end

       6005 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6005");
      end

       6006 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6006");
      end

       6007 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6007");
      end

       6008 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6008");
      end

       6009 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  6009");
      end

       6010 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6010");
      end

       6011 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6011");
      end

       6012 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6012");
      end

       6013 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6013");
      end

       6014 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6014");
      end

       6015 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6015");
      end

       6016 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6016");
      end

       6017 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6017");
      end

       6018 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6018");
      end

       6019 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6019");
      end

       6020 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6020");
      end

       6021 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6021");
      end

       6022 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  6022");
      end

       6023 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6023");
      end

       6024 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6024");
      end

       6025 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6025");
      end

       6026 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6026");
      end

       6027 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6027");
      end

       6028 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6028");
      end

       6029 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6029");
      end

       6030 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6030");
      end

       6031 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6031");
      end

       6032 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6032");
      end

       6033 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6033");
      end

       6034 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6034");
      end

       6035 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6035");
      end

       6036 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6036");
      end

       6037 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6037");
      end

       6038 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6038");
      end

       6039 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6039");
      end

       6040 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6040");
      end

       6041 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6041");
      end

       6042 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6042");
      end

       6043 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6043");
      end

       6044 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6044");
      end

       6045 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6045");
      end

       6046 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6046");
      end

       6047 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6047");
      end

       6048 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6048");
      end

       6049 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6049");
      end

       6050 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6050");
      end

       6051 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6051");
      end

       6052 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6052");
      end

       6053 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6053");
      end

       6054 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6054");
      end

       6055 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6055");
      end

       6056 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6056");
      end

       6057 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6057");
      end

       6058 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6058");
      end

       6059 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6059");
      end

       6060 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6060");
      end

       6061 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6061");
      end

       6062 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6062");
      end

       6063 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6063");
      end

       6064 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6064");
      end

       6065 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6065");
      end

       6066 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6066");
      end

       6067 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6067");
      end

       6068 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6068");
      end

       6069 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6069");
      end

       6070 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6070");
      end

       6071 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6071");
      end

       6072 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6072");
      end

       6073 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6073");
      end

       6074 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6074");
      end

       6075 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  6075");
      end

       6076 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6076");
      end

       6077 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6077");
      end

       6078 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6079;
      end

       6079 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2507] = localMem[2507] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6080;
      end

       6080 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 5582;
      end

       6081 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6081");
      end

       6082 :
      begin                                                                     // assert
if (0) begin
  $display("AAAA %4d %4d assert", steps, ip);
end
         $display("Should not be executed  6082");
      end

       6083 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6083");
      end

       6084 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6084");
      end

       6085 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6086;
      end

       6086 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2735] = heapMem[localMem[2376]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6087;
      end

       6087 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2736] = heapMem[localMem[2376]*7 + 1];
              updateArrayLength(2, 0, 0);
              ip = 6088;
      end

       6088 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2737] = heapMem[localMem[2376]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 6089;
      end

       6089 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2736] != 1 ? 6093 : 6090;
      end

       6090 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6090");
      end

       6091 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6091");
      end

       6092 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6092");
      end

       6093 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6094;
      end

       6094 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
              ip = localMem[2736] != 2 ? 6102 : 6095;
      end

       6095 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              localMem[2739] = localMem[2737] + 1;
              updateArrayLength(2, 0, 0);
              ip = 6096;
      end

       6096 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2740] = heapMem[localMem[2735]*7 + 4];
              updateArrayLength(2, 0, 0);
              ip = 6097;
      end

       6097 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2740] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2739], localMem[2740], arraySizes[localMem[2740]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2739] && i <= arraySizes[localMem[2740]]) begin
                  heapMem[NArea * localMem[2740] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2740] + localMem[2739]] = 6;                                    // Insert new value
              arraySizes[localMem[2740]] = arraySizes[localMem[2740]] + 1;                              // Increase array size
              ip = 6098;
      end

       6098 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2741] = heapMem[localMem[2735]*7 + 5];
              updateArrayLength(2, 0, 0);
              ip = 6099;
      end

       6099 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
//$display("AAAA %4d %4d shiftUp", steps, ip);
              for(i = 0; i < NArea; i = i + 1) arrayShift[i] = heapMem[NArea * localMem[2741] + i]; // Copy source array
//$display("BBBB pos=%d array=%d length=%d", localMem[2739], localMem[2741], arraySizes[localMem[2741]]);
              for(i = 0; i < NArea; i = i + 1) begin                            // Move original array up
                if (i > localMem[2739] && i <= arraySizes[localMem[2741]]) begin
                  heapMem[NArea * localMem[2741] + i] = arrayShift[i-1];
//$display("CCCC index=%d value=%d", i, arrayShift[i-1]);
                end
              end
              heapMem[NArea * localMem[2741] + localMem[2739]] = 66;                                    // Insert new value
              arraySizes[localMem[2741]] = arraySizes[localMem[2741]] + 1;                              // Increase array size
              ip = 6100;
      end

       6100 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[2735]*7 + 0] = heapMem[localMem[2735]*7 + 0] + 1;
              updateArrayLength(1, localMem[2735], 0);
              ip = 6101;
      end

       6101 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
              ip = 6108;
      end

       6102 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6102");
      end

       6103 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6103");
      end

       6104 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  6104");
      end

       6105 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6105");
      end

       6106 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  6106");
      end

       6107 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6107");
      end

       6108 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6109;
      end

       6109 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
              heapMem[localMem[0]*7 + 0] = heapMem[localMem[0]*7 + 0] + 1;
              updateArrayLength(1, localMem[0], 0);
              ip = 6110;
      end

       6110 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6111;
      end

       6111 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2745] = heapMem[localMem[2735]*7 + 0];
              updateArrayLength(2, 0, 0);
              ip = 6112;
      end

       6112 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2746] = heapMem[localMem[2735]*7 + 3];
              updateArrayLength(2, 0, 0);
              ip = 6113;
      end

       6113 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2747] = heapMem[localMem[2746]*7 + 2];
              updateArrayLength(2, 0, 0);
              ip = 6114;
      end

       6114 :
      begin                                                                     // jLt
if (0) begin
  $display("AAAA %4d %4d jLt", steps, ip);
end
              ip = localMem[2745] <  localMem[2747] ? 6334 : 6115;
      end

       6115 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6115");
      end

       6116 :
      begin                                                                     // shiftRight
if (0) begin
  $display("AAAA %4d %4d shiftRight", steps, ip);
end
         $display("Should not be executed  6116");
      end

       6117 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6117");
      end

       6118 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6118");
      end

       6119 :
      begin                                                                     // jEq
if (0) begin
  $display("AAAA %4d %4d jEq", steps, ip);
end
         $display("Should not be executed  6119");
      end

       6120 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6120");
      end

       6121 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6121");
      end

       6122 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6122");
      end

       6123 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6123");
      end

       6124 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6124");
      end

       6125 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6125");
      end

       6126 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6126");
      end

       6127 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6127");
      end

       6128 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6128");
      end

       6129 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6129");
      end

       6130 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6130");
      end

       6131 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  6131");
      end

       6132 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  6132");
      end

       6133 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6133");
      end

       6134 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6134");
      end

       6135 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6135");
      end

       6136 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6136");
      end

       6137 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6137");
      end

       6138 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6138");
      end

       6139 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6139");
      end

       6140 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6140");
      end

       6141 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6141");
      end

       6142 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6142");
      end

       6143 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6143");
      end

       6144 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6144");
      end

       6145 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6145");
      end

       6146 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6146");
      end

       6147 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6147");
      end

       6148 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6148");
      end

       6149 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6149");
      end

       6150 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6150");
      end

       6151 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  6151");
      end

       6152 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6152");
      end

       6153 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6153");
      end

       6154 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6154");
      end

       6155 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6155");
      end

       6156 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6156");
      end

       6157 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6157");
      end

       6158 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6158");
      end

       6159 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6159");
      end

       6160 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6160");
      end

       6161 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6161");
      end

       6162 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6162");
      end

       6163 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6163");
      end

       6164 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6164");
      end

       6165 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6165");
      end

       6166 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6166");
      end

       6167 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6167");
      end

       6168 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6168");
      end

       6169 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6169");
      end

       6170 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6170");
      end

       6171 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6171");
      end

       6172 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6172");
      end

       6173 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6173");
      end

       6174 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  6174");
      end

       6175 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6175");
      end

       6176 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6176");
      end

       6177 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6177");
      end

       6178 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6178");
      end

       6179 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6179");
      end

       6180 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6180");
      end

       6181 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6181");
      end

       6182 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6182");
      end

       6183 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6183");
      end

       6184 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6184");
      end

       6185 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6185");
      end

       6186 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6186");
      end

       6187 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6187");
      end

       6188 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6188");
      end

       6189 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6189");
      end

       6190 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6190");
      end

       6191 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6191");
      end

       6192 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6192");
      end

       6193 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6193");
      end

       6194 :
      begin                                                                     // assertNe
if (0) begin
  $display("AAAA %4d %4d assertNe", steps, ip);
end
         $display("Should not be executed  6194");
      end

       6195 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6195");
      end

       6196 :
      begin                                                                     // arrayIndex
if (0) begin
  $display("AAAA %4d %4d arrayIndex", steps, ip);
end
         $display("Should not be executed  6196");
      end

       6197 :
      begin                                                                     // subtract
if (0) begin
  $display("AAAA %4d %4d subtract", steps, ip);
end
         $display("Should not be executed  6197");
      end

       6198 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6198");
      end

       6199 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6199");
      end

       6200 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6200");
      end

       6201 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6201");
      end

       6202 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6202");
      end

       6203 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6203");
      end

       6204 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6204");
      end

       6205 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6205");
      end

       6206 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6206");
      end

       6207 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  6207");
      end

       6208 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6208");
      end

       6209 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  6209");
      end

       6210 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6210");
      end

       6211 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6211");
      end

       6212 :
      begin                                                                     // shiftUp
if (0) begin
  $display("AAAA %4d %4d shiftUp", steps, ip);
end
         $display("Should not be executed  6212");
      end

       6213 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6213");
      end

       6214 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6214");
      end

       6215 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6215");
      end

       6216 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6216");
      end

       6217 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6217");
      end

       6218 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6218");
      end

       6219 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6219");
      end

       6220 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6220");
      end

       6221 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6221");
      end

       6222 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6222");
      end

       6223 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6223");
      end

       6224 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6224");
      end

       6225 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6225");
      end

       6226 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6226");
      end

       6227 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6227");
      end

       6228 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6228");
      end

       6229 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6229");
      end

       6230 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6230");
      end

       6231 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6231");
      end

       6232 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6232");
      end

       6233 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6233");
      end

       6234 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6234");
      end

       6235 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6235");
      end

       6236 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6236");
      end

       6237 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6237");
      end

       6238 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6238");
      end

       6239 :
      begin                                                                     // not
if (0) begin
  $display("AAAA %4d %4d not", steps, ip);
end
         $display("Should not be executed  6239");
      end

       6240 :
      begin                                                                     // jNe
if (0) begin
  $display("AAAA %4d %4d jNe", steps, ip);
end
         $display("Should not be executed  6240");
      end

       6241 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6241");
      end

       6242 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6242");
      end

       6243 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6243");
      end

       6244 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6244");
      end

       6245 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6245");
      end

       6246 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6246");
      end

       6247 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6247");
      end

       6248 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6248");
      end

       6249 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6249");
      end

       6250 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6250");
      end

       6251 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6251");
      end

       6252 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6252");
      end

       6253 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6253");
      end

       6254 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6254");
      end

       6255 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6255");
      end

       6256 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6256");
      end

       6257 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6257");
      end

       6258 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6258");
      end

       6259 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6259");
      end

       6260 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6260");
      end

       6261 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6261");
      end

       6262 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6262");
      end

       6263 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6263");
      end

       6264 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6264");
      end

       6265 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6265");
      end

       6266 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6266");
      end

       6267 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6267");
      end

       6268 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6268");
      end

       6269 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6269");
      end

       6270 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6270");
      end

       6271 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  6271");
      end

       6272 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6272");
      end

       6273 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6273");
      end

       6274 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6274");
      end

       6275 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6275");
      end

       6276 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6276");
      end

       6277 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6277");
      end

       6278 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6278");
      end

       6279 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6279");
      end

       6280 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6280");
      end

       6281 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6281");
      end

       6282 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6282");
      end

       6283 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6283");
      end

       6284 :
      begin                                                                     // jGe
if (0) begin
  $display("AAAA %4d %4d jGe", steps, ip);
end
         $display("Should not be executed  6284");
      end

       6285 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6285");
      end

       6286 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6286");
      end

       6287 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6287");
      end

       6288 :
      begin                                                                     // add
if (0) begin
  $display("AAAA %4d %4d add", steps, ip);
end
         $display("Should not be executed  6288");
      end

       6289 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6289");
      end

       6290 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6290");
      end

       6291 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6291");
      end

       6292 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6292");
      end

       6293 :
      begin                                                                     // array
if (0) begin
  $display("AAAA %4d %4d array", steps, ip);
end
         $display("Should not be executed  6293");
      end

       6294 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6294");
      end

       6295 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6295");
      end

       6296 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6296");
      end

       6297 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6297");
      end

       6298 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6298");
      end

       6299 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6299");
      end

       6300 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6300");
      end

       6301 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6301");
      end

       6302 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6302");
      end

       6303 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6303");
      end

       6304 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6304");
      end

       6305 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6305");
      end

       6306 :
      begin                                                                     // moveLong
if (0) begin
  $display("AAAA %4d %4d moveLong", steps, ip);
end
         $display("Should not be executed  6306");
      end

       6307 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6307");
      end

       6308 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6308");
      end

       6309 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6309");
      end

       6310 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6310");
      end

       6311 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6311");
      end

       6312 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6312");
      end

       6313 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6313");
      end

       6314 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6314");
      end

       6315 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6315");
      end

       6316 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6316");
      end

       6317 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6317");
      end

       6318 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6318");
      end

       6319 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6319");
      end

       6320 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6320");
      end

       6321 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6321");
      end

       6322 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6322");
      end

       6323 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6323");
      end

       6324 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6324");
      end

       6325 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6325");
      end

       6326 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6326");
      end

       6327 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6327");
      end

       6328 :
      begin                                                                     // resize
if (0) begin
  $display("AAAA %4d %4d resize", steps, ip);
end
         $display("Should not be executed  6328");
      end

       6329 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6329");
      end

       6330 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6330");
      end

       6331 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
         $display("Should not be executed  6331");
      end

       6332 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
         $display("Should not be executed  6332");
      end

       6333 :
      begin                                                                     // jmp
if (0) begin
  $display("AAAA %4d %4d jmp", steps, ip);
end
         $display("Should not be executed  6333");
      end

       6334 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6335;
      end

       6335 :
      begin                                                                     // mov
if (0) begin
  $display("AAAA %4d %4d mov", steps, ip);
end
              localMem[2744] = 0;
              updateArrayLength(2, 0, 0);
              ip = 6336;
      end

       6336 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6337;
      end

       6337 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6338;
      end

       6338 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6339;
      end

       6339 :
      begin                                                                     // label
if (0) begin
  $display("AAAA %4d %4d label", steps, ip);
end
              ip = 6340;
      end

       6340 :
      begin                                                                     // free
if (0) begin
  $display("AAAA %4d %4d free", steps, ip);
end
                                 arraySizes[localMem[2376]] = 0;
              freedArrays[freedArraysTop] = localMem[2376];
              freedArraysTop = freedArraysTop + 1;
              ip = 6341;
      end
      default: begin
        success  = 1;
        finished = 1;
      end
    endcase
    if (steps <=    492) clock <= ~ clock;                                      // Must be non sequential to fire the next iteration
    if (0) begin
      for(i = 0; i < 200; i = i + 1) $write("%2d",   localMem[i]); $display("");
      for(i = 0; i < 200; i = i + 1) $write("%2d",    heapMem[i]); $display("");
      for(i = 0; i < 200; i = i + 1) $write("%2d", arraySizes[i]); $display("");
    end
  end
endmodule
