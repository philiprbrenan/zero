  parameter integer NInstructions = 4;

  task startTest();                                                             // Array_test: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000001101000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   2] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   3] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
    end
  endtask

  task endTest();                                                               // Array_test: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 11;
    end
  endtask
