  parameter integer NInstructions = 2;

  task startTest();                                                             // Subtract_test: load code
    begin

      code[   0] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000010000000000010000000000;                                          // subtract
      code[   1] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
    end
  endtask

  task endTest();                                                               // Subtract_test: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 2;
    end
  endtask
