  parameter integer NInstructions = 1141;

  task startTest();                                                             // BTree: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[   2] = 'b0000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // inSize
      code[   3] = 'b0000000000000000000000000001100000000000000000000000000000000000000000000000000000100000100011100000000011000000100001000000000000000000000000000000000000000000000000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jFalse
      code[   4] = 'b0000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000001000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // in
      code[   5] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000111000000000000000100000100001000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[   6] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100001000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   7] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110000000000000001000000101010000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   8] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110000000000000011000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   9] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110000000000000000000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  10] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110000000000000010000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  11] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000100000111001100000000001000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[  12] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  13] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000100000101110000000000010100000100001000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // jNe
      code[  14] = 'b0000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000000100000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // in
      code[  15] = 'b0000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000000000000010100000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // in
      code[  16] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  17] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  18] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011100000100001000000000000000000000000000000000011000000000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  19] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000110010000000000001010000100001000000000000000000000000000000000000000000000000001110000010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[  20] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  21] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000000000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  22] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  23] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010010000100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  24] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000000100000101010000000000000000000000000000000000000000000000000001001000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  25] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001010000100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  26] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000010100000101010000000000000000000000000000000000000000000000000000101000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  27] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  28] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000011000000101010000000000000000000000000000000000000000000000000001100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  29] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000010000000101010000000000000000000000000000000000011000000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  30] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000100000000000010000000101010000000000000000000000000000000000011000000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  31] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011010000100001000000000000000000000000000000000000010000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  32] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110100000000000000000000101010000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  33] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110000100001000000000000000000000000000000000000010000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  34] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001100000000000000000000101010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  35] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000101010000000000000000000000000000000000011000000000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  36] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110000000000000011000000101010000000000000000000000000000000000000000000000000000001000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  37] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000100000010000000000000010010000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[  38] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  39] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110000100001000000000000000000000000000000000011100000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  40] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110000100001000000000000000000000000000000000011000000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  41] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000100001000000000011010000100001000000000000000000000000000000000000000000000000001011000010000100000000000000000000000000000000000000000000000000011100001000010000000000;                                          // jGe
      code[  42] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110000100001000000000000000000000000000000000011100000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  43] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000011110000000000000110000100001000000000000000000000000000000000000000000000000001111000010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[  44] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000000001000100001000000000000000000000000000000000011100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[  45] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000110110000000000010110000100001000000000000000000000000000000000000000000000000000000100010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[  46] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001000100001000000000000000000000000000000000011100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  47] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000001001000100001000000000000000000000000000000000000000000000000001000100010000100000000000000000000000000000000000000000000000000001000001000010000000000;                                          // arrayIndex
      code[  48] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000001110000100001000000000000000000000000000000000000000000000000000100100010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[  49] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000001001000100001000000000000000000000000000000000000000000000000000100100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[  50] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011001000100001000000000000000000000000000000000011100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  51] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110010000000000001001000011010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  52] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000011000000110011110000000010010000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[  53] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  54] = 'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000101000100001000000000000000000000000000000000000000000000000001000100010000100000000000000000000000000000000000000000000000000001000001000010000000000;                                          // arrayCountGreater
      code[  55] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000100000000000011110000100001000000000000000000000000000000000000000000000000000010100010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[  56] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010101000100001000000000000000000000000000000000011100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  57] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010000000000010110000011010000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  58] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001101000100001000000000000000000000000000000000011100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  59] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011010000000000010110000011010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  60] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000101010000000000000000000000000000000000000000000000000001011000010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  61] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000101010000000000000000000000000000000000011000000000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  62] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000011000000100101110000000010010000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[  63] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  64] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000011101000100001000000000000000000000000000000000000000000000000001000100010000100000000000000000000000000000000000000000000000000001000001000010000000000;                                          // arrayCountLess
      code[  65] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000011000100001000000000000000000000000000000000011100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  66] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000110000000000011101000011010000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[  67] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010011000100001000000000000000000000000000000000011100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  68] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000100110000000000011101000011010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[  69] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000101010000000000000000000000000000000000011100000000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  70] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000101010000000000000000000000000000000000011000000000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  71] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000011000000000001110000000010010000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[  72] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  73] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  74] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  75] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011000100001000000000000000000000000000000000011000000000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  76] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  77] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000111000100001000000000000000000000000000000000001011000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  78] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111000100001000000000000000000000000000000000001011000000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  79] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111000100001000000000000000000000000000000000010111000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  80] = 'b0000000000000000000000000011100000000000000000000000000000000000000000000000000000000000001110110000000001001000100001000000000000000000000000000000000000000000000000000011100010000100000000000000000000000000000000000000000000000000011110001000010000000000;                                          // jLt
      code[  81] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111000100001000000000000000000000000000000000000000000000000000111100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  82] = 'b0000000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000000000000011111000100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftRight
      code[  83] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  84] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000100100001000000000000000000000000000000000001011000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  85] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000100001100000000000101000100001000000000000000000000000000000000000000000000000001000010010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[  86] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000100100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  87] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000000000000101010000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  88] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  89] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011000100100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  90] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000000100000101010000000000000000000000000000000000000000000000000001100010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  91] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100100100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[  92] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000010100000101010000000000000000000000000000000000000000000000000000010010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  93] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  94] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000011000000101010000000000000000000000000000000000000000000000000001011100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  95] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000000010000000101010000000000000000000000000000000000010111000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[  96] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000010000000101010000000000000000000000000000000000010111000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  97] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000010100100100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[  98] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000101110000000000010101000100001000000000000000000000000000000000000000000000000001010010010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[  99] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001100100100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 100] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000001100000101010000000000000000000000000000000000000000000000000000110010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 101] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011100100100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 102] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000010100100001000000000000000000000000000000000001000100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 103] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000101000000000000000000101010000000000000000000000000000000000011100100000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 104] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010010100100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 105] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001010100100001000000000000000000000000000000000001000100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 106] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000010101000000000000000000101010000000000000000000000000000000000010010100000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 107] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011010100100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 108] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110100100001000000000000000000000000000000000001000100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 109] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110100100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 110] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001101000000000000000000101010000000000000000000000000000000000011010100000000000000010001101000000000000000000000000000000000000000000000000000101101001000010000000000;                                          // moveLong
      code[ 111] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110100100001000000000000000000000000000000000001000100000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 112] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110100100001000000000000000000000000000000000000000000000000000111010010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 113] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000001100100001000000000000000000000000000000000001000100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 114] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 115] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001100100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 116] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 117] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000001011000100001000000000000000000000000000000000000000000000000001000110010000100000000000000000000000000000000000000000000000000111101001000010000000000;                                          // jGe
      code[ 118] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001001100100001000000000000000000000000000000000000001100000000001000110001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 119] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010011000000000001000000101010000000000000000000000000000000000000000000000000000100010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 120] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 121] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001100100001000000000000000000000000000000000000000000000000001000110010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 122] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000000011000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 123] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 124] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011001100100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 125] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000011001100100001000000000000000000000000000000000000000000000000000000010010000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 126] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000100000000000001101000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 127] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 128] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000101100100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 129] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010101100100001000000000000000000000000000000000001000100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 130] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000101011000000000000000000101010000000000000000000000000000000000000101100000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 131] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001101100100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 132] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011101100100001000000000000000000000000000000000001000100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 133] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000111011000000000000000000101010000000000000000000000000000000000001101100000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 134] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 135] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010110000000000000000000101010000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 136] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010001000000000001000000101010000000000000000000000000000000000000000000000000001000010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 137] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000011100100001000000000000000000000000000000000010000100000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 138] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010011100100001000000000000000000000000000000000010000100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 139] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011100100001000000000000000000000000000000000010011100000000000001110001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 140] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000110010000000000011011000100001000000000000000000000000000000000000000000000000000101110010000100000000000000000000000000000000000000000000000000010110001000010000000000;                                          // jNe
      code[ 141] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011100100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 142] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000111100100001000000000000000000000000000000000011011100000000001111100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 143] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111100100001000000000000000000000000000000000010000100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 144] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101111000000000000011100011010000000000000000000000000000000000000000000000000000011110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 145] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111100100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 146] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111100100001000000000000000000000000000000000001111100000000001111100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 147] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000010100001000000000000000000000000000000000010000100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 148] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000100000000000011100011010000000000000000000000000000000000000000000000000001111110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 149] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000010100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 150] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000010000010100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 151] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000010100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 152] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000001000010100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 153] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010100001000000000000000000000000000000000000000000000000000001110010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 154] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100001000000000000000000101010000000000000000000000000000000000000000000000000001100001010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 155] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000100010100001000000000000000000000000000000000010000100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 156] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000100000000011000010011010000000000000000000000000000000000000000000000000000100010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 157] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001100010000000010001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 158] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111010000000000000111000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 159] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 160] = 'b0000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000010010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // assertNe
      code[ 161] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010100010100001000000000000000000000000000000000010000100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 162] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000001100010100001000000000000000000000000000000000000000000000000001010001010000100000000000000000000000000000000000000000000000000010110001000010000000000;                                          // arrayIndex
      code[ 163] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000001100010100001000000000000000000000000000000000000000000000000000110001010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 164] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011100010100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 165] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000010010100001000000000000000000000000000000000011100010000000001111100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 166] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010010010100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 167] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001010010100001000000000000000000000000000000000010010010000000001111100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 168] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011010010100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 169] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000011010010100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 170] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110010100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 171] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000000110010100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 172] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110010100001000000000000000000000000000000000010000100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 173] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000101100100000000001100010011010000000000000000000000000000000000000000000000000000001001010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 174] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110010100001000000000000000000000000000000000010000100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 175] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000011100100000000001100010011010000000000000000000000000000000000000000000000000000101001010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 176] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110010100001000000000000000000000000000000000010000100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 177] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001000000000000000000000000000000000000000000000000000110001010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 178] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000111100100000000000001010011010000000000000000000000000000000000000000000000000000100010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 179] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000101010000000000000000000000000000000000010000100000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 180] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000101011100000000010001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 181] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 182] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 183] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010001010100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 184] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000000000000101010000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 185] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 186] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001001010100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 187] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000000100000101010000000000000000000000000000000000000000000000000000100101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 188] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011001010100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 189] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000010100000101010000000000000000000000000000000000000000000000000001100101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 190] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 191] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000011000000101010000000000000000000000000000000000000000000000000001011100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 192] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000000010000000101010000000000000000000000000000000000010111000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 193] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000010000000101010000000000000000000000000000000000010111000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 194] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 195] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000000000000101010000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 196] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 197] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 198] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000000100000101010000000000000000000000000000000000000000000000000001010101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 199] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001101010100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 200] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000010100000101010000000000000000000000000000000000000000000000000000110101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 201] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 202] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000011000000101010000000000000000000000000000000000000000000000000001011100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 203] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000000010000000101010000000000000000000000000000000000010111000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 204] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000010000000101010000000000000000000000000000000000010111000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 205] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000011101010100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 206] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000001011000000000010111000100001000000000000000000000000000000000000000000000000001110101010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 207] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000011010100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 208] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000001100000101010000000000000000000000000000000000000000000000000000001101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 209] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010011010100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 210] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000001100000101010000000000000000000000000000000000000000000000000001001101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 211] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011010100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 212] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011010100001000000000000000000000000000000000010001010000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 213] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000110110100000000000000000101010000000000000000000000000000000000001011010000000000000000010101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 214] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000111010100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 215] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111010100001000000000000000000000000000000000010001010000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 216] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000101110100000000000000000101010000000000000000000000000000000000000111010000000000000000010101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 217] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111010100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 218] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111010100001000000000000000000000000000000000010001010000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 219] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 220] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000111110100000000000000000101010000000000000000000000000000000000001111010000000000000000010101000000000000000000000000000000000000000000000000000000001101000010000000000;                                          // moveLong
      code[ 221] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000110100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 222] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000110100001000000000000000000000000000000000000101010000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 223] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000010001100000000000000000101010000000000000000000000000000000000010000110000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 224] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011000110100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 225] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000100110100001000000000000000000000000000000000000101010000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 226] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001100000000000000000101010000000000000000000000000000000000011000110000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 227] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010100110100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 228] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001100110100001000000000000000000000000000000000000101010000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 229] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100110100001000000000000000000000000000000000000000000000000001111100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 230] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000011001100000000000000000101010000000000000000000000000000000000010100110000000000000010001101000000000000000000000000000000000000000000000000000111001101000010000000000;                                          // moveLong
      code[ 231] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000010110100001000000000000000000000000000000000010001010000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 232] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010110100001000000000000000000000000000000000000000000000000000001011010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 233] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001010110100001000000000000000000000000000000000010001010000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 234] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 235] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011010110100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 236] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 237] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000001000100100001000000000000000000000000000000000000000000000000001101011010000100000000000000000000000000000000000000000000000000100101101000010000000000;                                          // jGe
      code[ 238] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110110100001000000000000000000000000000000000001010110000000001101011001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 239] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001101100000000001000000101010000000000000000000000000000000000000000000000000001000101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 240] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 241] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010110100001000000000000000000000000000000000000000000000000001101011010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 242] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000000000100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 243] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 244] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110110100001000000000000000000000000000000000000101010000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 245] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110110100001000000000000000000000000000000000000000000000000001011011010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 246] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110110100001000000000000000000000000000000000000101010000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 247] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 248] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000001110100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 249] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 250] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000001100100100001000000000000000000000000000000000000000000000000000000111010000100000000000000000000000000000000000000000000000000011101101000010000000000;                                          // jGe
      code[ 251] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001110100001000000000000000000000000000000000011110110000000000000111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 252] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100011100000000001000000101010000000000000000000000000000000000000000000000000000010101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 253] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 254] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100001000000000000000000000000000000000000000000000000000000111010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 255] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000000100100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 256] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 257] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000010000000000001111000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 258] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 259] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001001110100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 260] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010110000000000001100000101010000000000000000000000000000000000000000000000000000100111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 261] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011001110100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 262] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000101110100001000000000000000000000000000000000010001010000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 263] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001011100000000000000000101010000000000000000000000000000000000011001110000000000000000010101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 264] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010101110100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 265] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001101110100001000000000000000000000000000000000010001010000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 266] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000011011100000000000000000101010000000000000000000000000000000000010101110000000000000000010101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 267] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011101110100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 268] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000011110100001000000000000000000000000000000000000101010000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 269] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000111100000000000000000101010000000000000000000000000000000000011101110000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 270] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010011110100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 271] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011110100001000000000000000000000000000000000000101010000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 272] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000010111100000000000000000101010000000000000000000000000000000000010011110000000000000010001101000000000000000000000000000000000000000000000000000111110001000010000000000;                                          // moveLong
      code[ 273] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 274] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100010100000000001000000101010000000000000000000000000000000000000000000000000000101100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 275] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010100000000001000000101010000000000000000000000000000000000000000000000000000101100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 276] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011110100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 277] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000111110100001000000000000000000000000000000000011011110000000001111100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 278] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111110100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 279] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111110100001000000000000000000000000000000000010111110000000001111100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 280] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111110100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 281] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111111100000000000000000101010000000000000000000000000000000000000000000000000000011111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 282] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000001100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 283] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000010000000000000000101010000000000000000000000000000000000000000000000000000111111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 284] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000001100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 285] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100000010000000000000000101010000000000000000000000000000000000000000000000000001000101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 286] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000001100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 287] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010000010000000010000000101010000000000000000000000000000000000000000000000000000010101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 288] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010110000000000000000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 289] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011000001100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 290] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000011000001100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 291] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000100001100001000000000000000000000000000000000001011000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 292] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000000100001100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 293] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010100001100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 294] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000010100001100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 295] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000010000000000000010001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 296] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011000000000000011001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 297] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 298] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011000100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 299] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000011001000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 300] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 301] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011000100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 302] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 303] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 304] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 305] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001100001100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 306] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 307] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000010000000010011110000000001110100100001000000000000000000000000000000000000000000000000000110000110000100000000000000000000000000000000000000000000000000110001100000010000000000;                                          // jGe
      code[ 308] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011100001100001000000000000000000000000000000000001011000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 309] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000000010001100001000000000000000000000000000000000000000000000000001110000110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 310] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010010001100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 311] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001010001100001000000000000000000000000000000000010010001000000000001000101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 312] = 'b0000000000000000000000001101100000000000000000000000000000000000000000000000000000000000100011110000000011110100100001000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000010100011000010000000000;                                          // jLe
      code[ 313] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000011010001100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 314] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000000001100100001000000000000000000000000000000000000000000000000001101000110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[ 315] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000000000000101010000000000000000000000000000000000000000000000000000101100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 316] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000010000000101010000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 317] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000011000000000000001000000101010000000000000000000000000000000000000000000000000001110000110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 318] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000010000000110101110000000001010100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 319] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 320] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110001100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 321] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110001100001000000000000000000000000000000000000110001000000001110000101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 322] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 323] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110001100001000000000000000000000000000000000010110001000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 324] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000001001100001000000000000000000000000000000000010110001000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 325] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001001100001000000000000000000000000000000000000001001000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 326] = 'b0000000000000000000000000011100000000000000000000000000000000000000000000000000000000000001110110000000011001100100001000000000000000000000000000000000000000000000000001111000110000100000000000000000000000000000000000000000000000000100010011000010000000000;                                          // jLt
      code[ 327] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001001001100001000000000000000000000000000000000000000000000000001000100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 328] = 'b0000000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000000000000001001001100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftRight
      code[ 329] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 330] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000101001100001000000000000000000000000000000000010110001000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 331] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000100001100000000010101100100001000000000000000000000000000000000000000000000000000010100110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[ 332] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010101001100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 333] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000000000000101010000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 334] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 335] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001101001100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 336] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000000100000101010000000000000000000000000000000000000000000000000000110100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 337] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011101001100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 338] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000010100000101010000000000000000000000000000000000000000000000000001110100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 339] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 340] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000011000000101010000000000000000000000000000000000000000000000000000000100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 341] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000000101010000000000000000000000000000000000000001001000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 342] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000010000000101010000000000000000000000000000000000000001001000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 343] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000000011001100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 344] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000101110000000000001101100100001000000000000000000000000000000000000000000000000000001100110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 345] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010011001100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 346] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000001100000101010000000000000000000000000000000000000000000000000001001100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 347] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011001100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 348] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011001100001000000000000000000000000000000000010101001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 349] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000110110010000000000000000101010000000000000000000000000000000000001011001000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 350] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000111001100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 351] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111001100001000000000000000000000000000000000010101001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 352] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000101110010000000000000000101010000000000000000000000000000000000000111001000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 353] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111001100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 354] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111001100001000000000000000000000000000000000010101001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 355] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 356] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000111110010000000000000000101010000000000000000000000000000000000001111001000000001100100101101000000000000000000000000000000000000000000000000000000001011000010000000000;                                          // moveLong
      code[ 357] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000101100001000000000000000000000000000000000010101001000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 358] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101100001000000000000000000000000000000000000000000000000001000010110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 359] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011000101100001000000000000000000000000000000000010101001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 360] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 361] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000100101100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 362] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 363] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000011011100100001000000000000000000000000000000000000000000000000000010010110000100000000000000000000000000000000000000000000000000010001011000010000000000;                                          // jGe
      code[ 364] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010100101100001000000000000000000000000000000000011000101000000000010010101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 365] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101001010000000001000000101010000000000000000000000000000000000000000000000000001010100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 366] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 367] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101100001000000000000000000000000000000000000000000000000000010010110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 368] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000010011100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 369] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 370] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001100101100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 371] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000001100101100001000000000000000000000000000000000000000000000000001100100110000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 372] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000100000000000011101100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 373] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 374] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011100101100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 375] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000010101100001000000000000000000000000000000000010101001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 376] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000101010000000000000000101010000000000000000000000000000000000011100101000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 377] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010010101100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 378] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001010101100001000000000000000000000000000000000010101001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 379] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000010101010000000000000000101010000000000000000000000000000000000010010101000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 380] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 381] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101100010000000000000000101010000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 382] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101010010000000001000000101010000000000000000000000000000000000000000000000000000010100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 383] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011010101100001000000000000000000000000000000000000101001000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 384] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110101100001000000000000000000000000000000000000101001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 385] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110101100001000000000000000000000000000000000000110101000000001101010101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 386] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000110010000000000000111100100001000000000000000000000000000000000000000000000000001011010110000100000000000000000000000000000000000000000000000000101100011000010000000000;                                          // jNe
      code[ 387] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110101100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 388] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110101100001000000000000000000000000000000000001110101000000000100100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 389] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000001101100001000000000000000000000000000000000000101001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 390] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000011010000000011010101011010000000000000000000000000000000000000000000000000001111010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 391] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001101100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 392] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001001101100001000000000000000000000000000000000010001101000000000100100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 393] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011001101100001000000000000000000000000000000000000101001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 394] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110011010000000011010101011010000000000000000000000000000000000000000000000000000100110110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 395] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000101101100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 396] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000000101101100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 397] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010101101100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 398] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000010101101100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 399] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101101100001000000000000000000000000000000000000000000000000001101010110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 400] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001010010000000000000000101010000000000000000000000000000000000000000000000000000110110110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 401] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011101101100001000000000000000000000000000000000000101001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 402] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111011010000000001101101011010000000000000000000000000000000000000000000000000001010100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 403] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001100010000000001001100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 404] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111010000000000010111100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 405] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 406] = 'b0000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010100110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // assertNe
      code[ 407] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000011101100001000000000000000000000000000000000000101001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 408] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000010011101100001000000000000000000000000000000000000000000000000000001110110000100000000000000000000000000000000000000000000000000101100011000010000000000;                                          // arrayIndex
      code[ 409] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000010011101100001000000000000000000000000000000000000000000000000001001110110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 410] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011101100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 411] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011101100001000000000000000000000000000000000001011101000000000100100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 412] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000111101100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 413] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111101100001000000000000000000000000000000000000111101000000000100100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 414] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111101100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 415] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000001111101100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 416] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111101100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 417] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000011111101100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 418] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000011100001000000000000000000000000000000000000101001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 419] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000110000000010011101011010000000000000000000000000000000000000000000000000001101110110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 420] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000011100001000000000000000000000000000000000000101001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 421] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000100000110000000010011101011010000000000000000000000000000000000000000000000000001011110110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 422] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000011100001000000000000000000000000000000000000101001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 423] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011100001000000000000000000000000000000000000000000000000001001110110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 424] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000000000000010000110000000011000011011010000000000000000000000000000000000000000000000000001010100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 425] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010000000000000000101010000000000000000000000000000000000000101001000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 426] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000101011100000000001001100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 427] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 428] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 429] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100011100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 430] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000000000000101010000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 431] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 432] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010100011100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 433] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000000100000101010000000000000000000000000000000000000000000000000001010001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 434] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001100011100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 435] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000010100000101010000000000000000000000000000000000000000000000000000110001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 436] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 437] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000011000000101010000000000000000000000000000000000000000000000000000000100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 438] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000000101010000000000000000000000000000000000000001001000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 439] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000010000000101010000000000000000000000000000000000000001001000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 440] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 441] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000000000000101010000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 442] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 443] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010011100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 444] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000000100000101010000000000000000000000000000000000000000000000000000001001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 445] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010010011100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 446] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000010100000101010000000000000000000000000000000000000000000000000001001001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 447] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 448] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000011000000101010000000000000000000000000000000000000000000000000000000100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 449] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000000101010000000000000000000000000000000000000001001000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 450] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000010000000101010000000000000000000000000000000000000001001000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 451] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000001010011100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 452] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000001011000000000001111100100001000000000000000000000000000000000000000000000000000101001110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 453] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000011010011100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 454] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000001100000101010000000000000000000000000000000000000000000000000001101001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 455] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000110011100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 456] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000001100000101010000000000000000000000000000000000000000000000000000011001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 457] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110011100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 458] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110011100001000000000000000000000000000000000000100011000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 459] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000011100110000000000000000101010000000000000000000000000000000000010110011000000000000000010101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 460] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110011100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 461] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000001011100001000000000000000000000000000000000000100011000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 462] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000010110000000000000000101010000000000000000000000000000000000011110011000000000000000010101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 463] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001011100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 464] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001001011100001000000000000000000000000000000000000100011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 465] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001011100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 466] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000010010110000000000000000101010000000000000000000000000000000000010001011000000000000000010101000000000000000000000000000000000000000000000000000110010111000010000000000;                                          // moveLong
      code[ 467] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000101011100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 468] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010101011100001000000000000000000000000000000000011100011000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 469] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000101010110000000000000000101010000000000000000000000000000000000000101011000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 470] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001101011100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 471] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011101011100001000000000000000000000000000000000011100011000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 472] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000111010110000000000000000101010000000000000000000000000000000000001101011000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 473] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000011011100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 474] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010011011100001000000000000000000000000000000000011100011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 475] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011100001000000000000000000000000000000000000000000000000000100100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 476] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000100110110000000000000000101010000000000000000000000000000000000000011011000000001100100101101000000000000000000000000000000000000000000000000000010110111000010000000000;                                          // moveLong
      code[ 477] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011011011100001000000000000000000000000000000000000100011000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 478] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011100001000000000000000000000000000000000000000000000000001101101110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 479] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111011100001000000000000000000000000000000000000100011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 480] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 481] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111011100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 482] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 483] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000011000010100001000000000000000000000000000000000000000000000000000111101110000100000000000000000000000000000000000000000000000000001110111000010000000000;                                          // jGe
      code[ 484] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111011100001000000000000000000000000000000000010111011000000000111101101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 485] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111110110000000001000000101010000000000000000000000000000000000000000000000000000010001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 486] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 487] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011100001000000000000000000000000000000000000000000000000000111101110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 488] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000010000010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 489] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 490] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000111100001000000000000000000000000000000000011100011000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 491] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111100001000000000000000000000000000000000000000000000000000000011110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 492] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000111100001000000000000000000000000000000000011100011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 493] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 494] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011000111100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 495] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 496] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000011100010100001000000000000000000000000000000000000000000000000001100011110000100000000000000000000000000000000000000000000000000100001111000010000000000;                                          // jGe
      code[ 497] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000100111100001000000000000000000000000000000000001000111000000001100011101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 498] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001001110000000001000000101010000000000000000000000000000000000000000000000000001110001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 499] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 500] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000111100001000000000000000000000000000000000000000000000000001100011110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 501] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000010100010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 502] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 503] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000010000000000011111100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 504] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 505] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010100111100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 506] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101100010000000001100000101010000000000000000000000000000000000000000000000000001010011110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 507] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001100111100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 508] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011100111100001000000000000000000000000000000000000100011000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 509] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000111001110000000000000000101010000000000000000000000000000000000001100111000000000000000010101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 510] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000010111100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 511] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010010111100001000000000000000000000000000000000000100011000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 512] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000100101110000000000000000101010000000000000000000000000000000000000010111000000000000000010101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 513] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001010111100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 514] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011010111100001000000000000000000000000000000000011100011000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 515] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000110101110000000000000000101010000000000000000000000000000000000001010111000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 516] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000110111100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 517] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010110111100001000000000000000000000000000000000011100011000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 518] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000101101110000000000000000101010000000000000000000000000000000000000110111000000001100100101101000000000000000000000000000000000000000000000000000010010011000010000000000;                                          // moveLong
      code[ 519] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 520] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001000110000000001000000101010000000000000000000000000000000000000000000000000001011000110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 521] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000111000110000000001000000101010000000000000000000000000000000000000000000000000001011000110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 522] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110111100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 523] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011110111100001000000000000000000000000000000000001110111000000000100100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 524] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000001111100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 525] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010001111100001000000000000000000000000000000000000001111000000000100100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 526] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001001111100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 527] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000010011110000000000000000101010000000000000000000000000000000000000000000000000001111011110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 528] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011001111100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 529] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000110011110000000000000000101010000000000000000000000000000000000000000000000000001000111110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 530] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000101111100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 531] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000001011110000000000000000101010000000000000000000000000000000000000000000000000000010001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 532] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010101111100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 533] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101011110000000010000000101010000000000000000000000000000000000000000000000000001110001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 534] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000101100010000000000000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 535] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001101111100001000000000000000000000000000000000010110001000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 536] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000001101111100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 537] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011101111100001000000000000000000000000000000000010110001000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 538] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000011101111100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 539] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000011111100001000000000000000000000000000000000010110001000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 540] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000000011111100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 541] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000010000000000000001001100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 542] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011000000000000000101100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 543] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 544] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110001100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 545] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000000101100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 546] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 547] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001110001100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 548] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 549] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000010000000000000000010010100001000000000000000000000000000000000000000000000000000111000110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 550] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011000100001000000000000000000000000000000000000000000000000001011000110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 551] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 552] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000010111110000000010110100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 553] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 554] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010011111100001000000000000000000000000000000000001011000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 555] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000001011111100001000000000000000000000000000000000000000000000000001001111110000100000000000000000000000000000000000000000000000000001000001000010000000000;                                          // arrayIndex
      code[ 556] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000010010010100001000000000000000000000000000000000000000000000000000101111110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[ 557] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000000000000101010000000000000000000000000000000000000000000000000000101100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 558] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000010000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 559] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000011000000000000001000000101010000000000000000000000000000000000000000000000000000101111110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 560] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000100111110000000001010100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 561] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 562] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000011011111100001000000000000000000000000000000000000000000000000001001111110000100000000000000000000000000000000000000000000000000001000001000010000000000;                                          // arrayCountLess
      code[ 563] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000000111111100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 564] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000001010010100001000000000000000000000000000000000000000000000000000011111110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[ 565] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000000000000101010000000000000000000000000000000000000000000000000000101100010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 566] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000010000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 567] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011000000000000001000000101010000000000000000000000000000000000000000000000000001101111110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 568] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000100011110000000001010100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 569] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 570] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010111111100001000000000000000000000000000000000001011000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 571] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001111111100001000000000000000000000000000000000010111111000000001101111101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 572] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 573] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000000100001000000000000000000000000000000000001111111000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 574] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010000000100001000000000000000000000000000000000001111111000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 575] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000000100001000000000000000000000000001000000010000000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 576] = 'b0000000000000000000000000011100000000000000000000000000000000000000000000000000000000000001110110000000010110010100001000000000000000000000000000000000000000000100000000000000010000100000000000000000000000000000000000000000010000000010000001000010000000000;                                          // jLt
      code[ 577] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000000100001000000000000000000000000000000000000000000100000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 578] = 'b0000000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000001000000011000000100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftRight
      code[ 579] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 580] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100000100001000000000000000000000000000000000001111111000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 581] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000100001100000000011110010100001000000000000000000000000000000000000000000100000001010000010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[ 582] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001100000100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 583] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000000000000101010000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 584] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 585] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000011100000100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 586] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000000100000101010000000000000000000000000000000000000000000100000001110000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 587] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000010000100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 588] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000010100000101010000000000000000000000000000000000000000000100000000001000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 589] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 590] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000011000000101010000000000000000000000000000000000000000000100000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 591] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000010000000101010000000000000000000000000001000000010000000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 592] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000010000000101010000000000000000000000000001000000010000000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 593] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000001000000010010000100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 594] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000101110000000000000001010100001000000000000000000000000000000000000000000100000001001000010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 595] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001010000100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 596] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000001100000101010000000000000000000000000000000000000000000100000000101000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 597] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011010000100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 598] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110000100001000000000000000000000000001000000001100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 599] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000001100000000000000000000101010000000000000000000000000001000000011010000100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 600] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010110000100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 601] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001110000100001000000000000000000000000001000000001100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 602] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000011100000000000000000000101010000000000000000000000000001000000010110000100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 603] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110000100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 604] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001000100001000000000000000000000000001000000001100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 605] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001000100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 606] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000000010000000000000000000101010000000000000000000000000001000000011110000100000000010000001101000000000000000000000000000000000000000000010000000100010001000010000000000;                                          // moveLong
      code[ 607] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001001000100001000000000000000000000000001000000001100000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 608] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011001000100001000000000000000000000000000000000000000000100000000100100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 609] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000101000100001000000000000000000000000001000000001100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 610] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 611] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010101000100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 612] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 613] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000010101010100001000000000000000000000000000000000000000000100000001010100010000100000000000000000000000000000000000000000010000000110010001000010000000000;                                          // jGe
      code[ 614] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001101000100001000000000000000000000000001000000000101000100000001010100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 615] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011010000000000001000000101010000000000000000000000000000000000000000000100000000110000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 616] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 617] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101000100001000000000000000000000000000000000000000000100000001010100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 618] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000011001010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 619] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 620] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011101000100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 621] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000011101000100001000000000000000000000000000000000000000000100000000010000010000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 622] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000100000000000010001010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 623] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 624] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000011000100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 625] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010011000100001000000000000000000000000001000000001100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 626] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000100110000000000000000000101010000000000000000000000000001000000000011000100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 627] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001011000100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 628] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011011000100001000000000000000000000000001000000001100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 629] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000110110000000000000000000101010000000000000000000000000001000000001011000100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 630] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 631] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011111110000000000000000101010000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 632] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011000000000000001000000101010000000000000000000000000000000000000000000100000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 633] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000111000100001000000000000000000000000001000000010100000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 634] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010111000100001000000000000000000000000001000000010100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 635] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001111000100001000000000000000000000000001000000010111000100000000011100001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 636] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000110010000000000001101010100001000000000000000000000000000000000000000000100000000111100010000100000000000000000000000000000000000000000000000000011111111000010000000000;                                          // jNe
      code[ 637] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111000100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 638] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000100100001000000000000000000000000001000000011111000100000001100000001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 639] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010000100100001000000000000000000000000001000000010100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 640] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100001001000000000111000011010000000000000000000000000000000000000000000100000000000010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 641] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000100100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 642] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000100100001000000000000000000000000001000000001000100100000001100000001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 643] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000100100100001000000000000000000000000001000000010100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 644] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001001001000000000111000011010000000000000000000000000000000000000000000100000001100010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 645] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100100100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 646] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000010100100100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 647] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001100100100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 648] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000001100100100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 649] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011100100100001000000000000000000000000000000000000000000100000000011100010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 650] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101000000000000000000000101010000000000000000000000000000000000000000000100000001110010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 651] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000010100100001000000000000000000000000001000000010100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 652] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000101001000000011100100011010000000000000000000000000000000000000000000100000000110000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 653] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001100010000000000110010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 654] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111010000000000011101010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 655] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 656] = 'b0000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000001010000010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // assertNe
      code[ 657] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010010100100001000000000000000000000000001000000010100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 658] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000001000000001010100100001000000000000000000000000000000000000000000100000001001010010000100000000000000000000000000000000000000000000000000011111111000010000000000;                                          // arrayIndex
      code[ 659] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000001000000001010100100001000000000000000000000000000000000000000000100000000101010010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 660] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011010100100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 661] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110100100001000000000000000000000000001000000011010100100000001100000001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 662] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010110100100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 663] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001110100100001000000000000000000000000001000000010110100100000001100000001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 664] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110100100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 665] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000011110100100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 666] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001100100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 667] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000000001100100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 668] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010001100100001000000000000000000000000001000000010100000000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 669] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000100011001000000001010100011010000000000000000000000000000000000000000000100000000011010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 670] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001001100100001000000000000000000000000001000000010100000000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 671] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000010011001000000001010100011010000000000000000000000000000000000000000000100000000111010010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 672] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001100100001000000000000000000000000001000000010100000000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 673] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101100100001000000000000000000000000000000000000000000100000000101010010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 674] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000110011001000000000101100011010000000000000000000000000000000000000000000100000000110000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 675] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000000000000000000000101010000000000000000000000000001000000010100000000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 676] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000101011100000000000110010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 677] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 678] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 679] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010101100100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 680] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000000000000101010000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 681] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 682] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001101100100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 683] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000000100000101010000000000000000000000000000000000000000000100000000110110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 684] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000011101100100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 685] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000010100000101010000000000000000000000000000000000000000000100000001110110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 686] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 687] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000011000000101010000000000000000000000000000000000000000000100000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 688] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000010000000101010000000000000000000000000001000000010000000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 689] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000010000000101010000000000000000000000000001000000010000000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 690] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000011100100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 691] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000000000000101010000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 692] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 693] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010011100100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 694] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000000100000101010000000000000000000000000000000000000000000100000001001110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 695] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001011100100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 696] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000010100000101010000000000000000000000000000000000000000000100000000101110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 697] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 698] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000011000000101010000000000000000000000000000000000000000000100000001000000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 699] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000010000000101010000000000000000000000000001000000010000000000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 700] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000010000000101010000000000000000000000000001000000010000000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 701] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000001000000011011100100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 702] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000001011000000000000011010100001000000000000000000000000000000000000000000100000001101110010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 703] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000111100100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 704] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000001100000101010000000000000000000000000000000000000000000100000000011110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 705] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010111100100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 706] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000001100000101010000000000000000000000000000000000000000000100000001011110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 707] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001111100100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 708] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111100100001000000000000000000000000001000000010101100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 709] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000111111000000000000000000101010000000000000000000000000001000000001111100000000000000000010101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 710] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000010100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 711] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010000010100001000000000000000000000000001000000010101100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 712] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000100000100000000000000000101010000000000000000000000000001000000000000010000000000000000010101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 713] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000010100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 714] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000010100001000000000000000000000000001000000010101100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 715] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100010100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 716] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000110000100000000000000000101010000000000000000000000000001000000001000010000000000000000010101000000000000000000000000000000000000000000010000000001000101000010000000000;                                          // moveLong
      code[ 717] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100010100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 718] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001100010100001000000000000000000000000001000000000011100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 719] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000011000100000000000000000101010000000000000000000000000001000000010100010100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 720] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011100010100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 721] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000010010100001000000000000000000000000001000000000011100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 722] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000000100100000000000000000101010000000000000000000000000001000000011100010100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 723] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010010010100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 724] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001010010100001000000000000000000000000001000000000011100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 725] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011010010100001000000000000000000000000000000000000000000100000001100000010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 726] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000010100100000000000000000101010000000000000000000000000001000000010010010100000000010000001101000000000000000000000000000000000000000000010000000110100101000010000000000;                                          // moveLong
      code[ 727] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110010100001000000000000000000000000001000000010101100000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 728] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010110010100001000000000000000000000000000000000000000000100000000011001010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 729] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001110010100001000000000000000000000000001000000010101100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 730] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 731] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110010100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 732] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 733] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000010111010100001000000000000000000000000000000000000000000100000001111001010000100000000000000000000000000000000000000000010000000101100101000010000000000;                                          // jGe
      code[ 734] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001010100001000000000000000000000000001000000001110010100000001111001001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 735] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000010100000000001000000101010000000000000000000000000000000000000000000100000001010110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 736] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 737] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011110010100001000000000000000000000000000000000000000000100000001111001010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 738] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000011011010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 739] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 740] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010001010100001000000000000000000000000001000000000011100000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 741] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001001010100001000000000000000000000000000000000000000000100000001000101010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 742] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001010100001000000000000000000000000001000000000011100000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 743] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 744] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000101010100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 745] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 746] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000010000110100001000000000000000000000000000000000000000000100000000010101010000100000000000000000000000000000000000000000010000000010010101000010000000000;                                          // jGe
      code[ 747] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010101010100001000000000000000000000000001000000011001010100000000010101001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 748] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101010100000000001000000101010000000000000000000000000000000000000000000100000000001110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 749] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 750] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101010100001000000000000000000000000000000000000000000100000000010101010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 751] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000011111010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 752] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 753] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000010000000000010011010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 754] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 755] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001101010100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 756] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011111110000000001100000101010000000000000000000000000000000000000000000100000000110101010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 757] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011101010100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 758] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000011010100001000000000000000000000000001000000010101100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 759] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000000110100000000000000000101010000000000000000000000000001000000011101010000000000000000010101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 760] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010011010100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 761] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001011010100001000000000000000000000000001000000010101100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 762] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000010110100000000000000000101010000000000000000000000000001000000010011010000000000000000010101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 763] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011011010100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 764] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000111010100001000000000000000000000000001000000000011100000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 765] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000001110100000000000000000101010000000000000000000000000001000000011011010100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 766] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010111010100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 767] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001111010100001000000000000000000000000001000000000011100000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 768] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000011110100000000000000000101010000000000000000000000000001000000010111010100000000010000001101000000000000000000000000000000000000000000010000000110000001000010000000000;                                          // moveLong
      code[ 769] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 770] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101011000000000001000000101010000000000000000000000000000000000000000000000000000111111110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 771] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000111000000000001000000101010000000000000000000000000000000000000000000000000000111111110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 772] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111010100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 773] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000110100001000000000000000000000000001000000011111010100000001100000001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 774] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010000110100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 775] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000110100001000000000000000000000000001000000010000110100000001100000001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 776] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000110100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 777] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000110001100000000000000000101010000000000000000000000000000000000000000000100000000000011010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 778] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000100110100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 779] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001001100000000000000000101010000000000000000000000000000000000000000000100000000100011010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 780] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100110100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 781] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101001100000000000000000101010000000000000000000000000000000000000000000100000001010110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 782] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001100110100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 783] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000011001100000000010000000101010000000000000000000000000000000000000000000100000000001110010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 784] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000011111110000000000000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 785] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011100110100001000000000000000000000000000000000001111111000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 786] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000011100110100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 787] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000010110100001000000000000000000000000000000000001111111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 788] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000000010110100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 789] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010010110100001000000000000000000000000000000000001111111000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 790] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000010010110100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 791] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000010000000000000000110010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 792] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011000000000000001110010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 793] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 794] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111111100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 795] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000001110010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 796] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 797] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011111111100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 798] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 799] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000010000000000000001000110100001000000000000000000000000000000000000000000000000001111111110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 800] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001011000100001000000000000000000000000000000000000000000000000000111111110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 801] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 802] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 803] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001100001000000000000000000000000000000000000000000000000000110000110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 804] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111101111111011100000000000000110100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 805] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 806] = 'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // assert
      code[ 807] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 808] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 809] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 810] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001010110100001000000000000000000000000000000000001100000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 811] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011010110100001000000000000000000000000000000000001100000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 812] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110110100001000000000000000000000000000000000001100000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 813] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000001000000000000011000110100001000000000000000000000000000000000000000000100000001101011010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // jNe
      code[ 814] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010110110100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 815] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101101101000000000110110011010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 816] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111011110000000010010000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 817] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 818] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000100000000000000100110100001000000000000000000000000000000000000000000100000001101011010000100000000000000000000000000000000000000000000000000010000000000010000000000;                                          // jNe
      code[ 819] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001110110100001000000000000000000000000000000000000000000100000000011011010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 820] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110110100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 821] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000111101101000000001110110011010000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 822] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001110100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 823] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000000011101000000001110110011010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 824] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010101100000000000000000101010000000000000000000000000001000000001010110000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 825] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111000000000000010100110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 826] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 827] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010001110100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 828] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000100011101000000000110110011010000000000000000000000000000000000000000000000000000010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 829] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001001110100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 830] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000010011101000000000110110011010000000000000000000000000000000000000000000000000001010000010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 831] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010101100000000000000000101010000000000000000000000000001000000001010110000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 832] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 833] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000101010000000000000000000000000000000000011000000000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 834] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 835] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000101110100001000000000000000000000000001000000001010110000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 836] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010101110100001000000000000000000000000001000000001010110000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 837] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001101110100001000000000000000000000000001000000010101110000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 838] = 'b0000000000000000000000000011100000000000000000000000000000000000000000000000000000000000001110110000000000010110100001000000000000000000000000000000000000000000100000000010111010000100000000000000000000000000000000000000000010000000011011101000010000000000;                                          // jLt
      code[ 839] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011101110100001000000000000000000000000000000000000000000100000000110111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 840] = 'b0000000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000001000000011101110100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftRight
      code[ 841] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000011110100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 842] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010011110100001000000000000000000000000001000000001010110000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 843] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000100001100000000001010110100001000000000000000000000000000000000000000000100000001001111010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[ 844] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001011110100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 845] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000000000000101010000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 846] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 847] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000011011110100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 848] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000000100000101010000000000000000000000000000000000000000000100000001101111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 849] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000111110100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 850] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000010100000101010000000000000000000000000000000000000000000100000000011111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 851] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 852] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000011000000101010000000000000000000000000000000000000000000100000001010111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 853] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101011100000000010000000101010000000000000000000000000001000000010101110000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 854] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000010000000101010000000000000000000000000001000000010101110000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 855] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000001000000010111110100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 856] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000101110000000000011010110100001000000000000000000000000000000000000000000100000001011111010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 857] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001111110100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 858] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000001100000101010000000000000000000000000000000000000000000100000000111111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 859] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111110100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 860] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000001100001000000000000000000000000001000000001011110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 861] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000000000010000000000000000101010000000000000000000000000001000000011111110100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 862] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010000001100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 863] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000001100001000000000000000000000000001000000001011110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 864] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000010000010000000000000000101010000000000000000000000000001000000010000001100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 865] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000001100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 866] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000100001100001000000000000000000000000001000000001011110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 867] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100001100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 868] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000001000010000000000000000101010000000000000000000000000001000000011000001100000000001111001101000000000000000000000000000000000000000000010000000101000011000010000000000;                                          // moveLong
      code[ 869] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001100001100001000000000000000000000000001000000001011110000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 870] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011100001100001000000000000000000000000000000000000000000100000000110000110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 871] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000010001100001000000000000000000000000001000000001011110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 872] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 873] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010010001100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 874] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 875] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000000001110100001000000000000000000000000000000000000000000100000001001000110000100000000000000000000000000000000000000000010000000111000011000010000000000;                                          // jGe
      code[ 876] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001010001100001000000000000000000000000001000000000010001100000001001000101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 877] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010100010000000001000000101010000000000000000000000000000000000000000000100000000101111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 878] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 879] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010010001100001000000000000000000000000000000000000000000100000001001000110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 880] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000001110110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 881] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 882] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011010001100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 883] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000011010001100001000000000000000000000000000000000000000000100000000001111010000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[ 884] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000100000000000000110110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 885] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 886] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110001100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 887] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010110001100001000000000000000000000000001000000001011110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 888] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000101100010000000000000000101010000000000000000000000000001000000000110001100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 889] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001110001100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 890] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110001100001000000000000000000000000001000000001011110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 891] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000111100010000000000000000101010000000000000000000000000001000000001110001100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 892] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 893] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010101100000000000000000101010000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 894] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010111100000000001000000101010000000000000000000000000000000000000000000100000001001111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 895] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001001100001000000000000000000000000001000000010011110000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 896] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010001001100001000000000000000000000000001000000010011110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 897] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001001001100001000000000000000000000000001000000010001001100000000000100101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 898] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000110010000000000010001110100001000000000000000000000000000000000000000000100000000100100110000100000000000000000000000000000000000000000010000000010101101000010000000000;                                          // jNe
      code[ 899] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001001100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 900] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000101001100001000000000000000000000000001000000011001001100000001110111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 901] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010101001100001000000000000000000000000001000000010011110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 902] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000101010011000000000001001011010000000000000000000000000000000000000000000100000000010100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 903] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001101001100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 904] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011101001100001000000000000000000000000001000000001101001100000001110111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 905] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000011001100001000000000000000000000000001000000010011110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 906] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000110011000000000001001011010000000000000000000000000000000000000000000100000001110100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 907] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010011001100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 908] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000010011001100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 909] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001011001100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 910] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000001011001100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 911] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011011001100001000000000000000000000000000000000000000000100000000000100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 912] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100111100000000000000000101010000000000000000000000000000000000000000000100000001101100110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 913] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000111001100001000000000000000000000000001000000010011110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 914] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001110011000000011011001011010000000000000000000000000000000000000000000100000000101111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 915] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001100010000000011100110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 916] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111010000000000001001110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 917] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 918] = 'b0000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000001001111010000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // assertNe
      code[ 919] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010111001100001000000000000000000000000001000000010011110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 920] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000001000000001111001100001000000000000000000000000000000000000000000100000001011100110000100000000000000000000000000000000000000000010000000010101101000010000000000;                                          // arrayIndex
      code[ 921] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000001000000001111001100001000000000000000000000000000000000000000000100000000111100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[ 922] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111001100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 923] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000101100001000000000000000000000000001000000011111001100000001110111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 924] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010000101100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 925] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000101100001000000000000000000000000001000000010000101100000001110111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 926] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000101100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 927] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000011000101100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[ 928] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000100101100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 929] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000000100101100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[ 930] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100101100001000000000000000000000000001000000010011110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 931] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000101001011000000001111001011010000000000000000000000000000000000000000000100000000000010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 932] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001100101100001000000000000000000000000001000000010011110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 933] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000011001011000000001111001011010000000000000000000000000000000000000000000100000000100010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 934] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011100101100001000000000000000000000000001000000010011110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 935] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010101100001000000000000000000000000000000000000000000100000000111100110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 936] = 'b0000000000000000000000000001110000000000000000000000000000000000000000000000000010000000111001011000000000010101011010000000000000000000000000000000000000000000100000000101111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // shiftUp
      code[ 937] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100111100000000000000000101010000000000000000000000000001000000010011110000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 938] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000101011100000000011100110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[ 939] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 940] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 941] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010010101100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 942] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000000000000101010000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 943] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 944] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001010101100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 945] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000000100000101010000000000000000000000000000000000000000000100000000101010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 946] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000011010101100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 947] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000010100000101010000000000000000000000000000000000000000000100000001101010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 948] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 949] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000011000000101010000000000000000000000000000000000000000000100000001010111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 950] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101011100000000010000000101010000000000000000000000000001000000010101110000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 951] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000010000000101010000000000000000000000000001000000010101110000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 952] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000110101100001000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 953] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000000000000101010000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 954] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 955] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010110101100001000000000000000000000000000000000000000000000000000110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 956] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000000100000101010000000000000000000000000000000000000000000100000001011010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 957] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001110101100001000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 958] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000010100000101010000000000000000000000000000000000000000000100000000111010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 959] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000001100000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 960] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000011000000101010000000000000000000000000000000000000000000100000001010111010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 961] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101011100000000010000000101010000000000000000000000000001000000010101110000000001000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 962] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000010000000101010000000000000000000000000001000000010101110000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 963] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000001000000011110101100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[ 964] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000001011000000000011001110100001000000000000000000000000000000000000000000100000001111010110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[ 965] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000001101100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 966] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000001100000101010000000000000000000000000000000000000000000100000000000110110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 967] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010001101100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[ 968] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000001100000101010000000000000000000000000000000000000000000100000001000110110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 969] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001001101100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 970] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001101100001000000000000000000000000001000000010010101000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 971] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000110011010000000000000000101010000000000000000000000000001000000001001101000000000000000010101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 972] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000101101100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 973] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010101101100001000000000000000000000000001000000010010101000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 974] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000101011010000000000000000101010000000000000000000000000001000000000101101000000000000000010101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 975] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001101101100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 976] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011101101100001000000000000000000000000001000000010010101000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 977] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000011101100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 978] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000111011010000000000000000101010000000000000000000000000001000000001101101000000000000000010101000000000000000000000000000000000000000000010000000000111011000010000000000;                                          // moveLong
      code[ 979] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010011101100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 980] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001011101100001000000000000000000000000001000000000110101000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 981] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000010111010000000000000000101010000000000000000000000000001000000010011101100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 982] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011011101100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 983] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000111101100001000000000000000000000000001000000000110101000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 984] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000001111010000000000000000101010000000000000000000000000001000000011011101100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[ 985] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010111101100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 986] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001111101100001000000000000000000000000001000000000110101000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 987] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011111101100001000000000000000000000000000000000000000000100000001110111010000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 988] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000011111010000000000000000101010000000000000000000000000001000000010111101100000000001111001101000000000000000000000000000000000000000000010000000111111011000010000000000;                                          // moveLong
      code[ 989] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000011100001000000000000000000000000001000000010010101000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 990] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000011100001000000000000000000000000000000000000000000100000000000001110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[ 991] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000011100001000000000000000000000000001000000010010101000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 992] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 993] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011000011100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 994] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 995] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000000011110100001000000000000000000000000000000000000000000100000001100001110000100000000000000000000000000000000000000000010000000100000111000010000000000;                                          // jGe
      code[ 996] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000100011100001000000000000000000000000001000000001000011100000001100001101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 997] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001000110000000001000000101010000000000000000000000000000000000000000000100000001001010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[ 998] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[ 999] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011000011100001000000000000000000000000000000000000000000100000001100001110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[1000] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000001101110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1001] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1002] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100011100001000000000000000000000000001000000000110101000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1003] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001100011100001000000000000000000000000000000000000000000100000001010001110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[1004] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011100011100001000000000000000000000000001000000000110101000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1005] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1006] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000010011100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1007] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1008] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011000000000000000111110100001000000000000000000000000000000000000000000100000000001001110000100000000000000000000000000000000000000000010000000011000111000010000000000;                                          // jGe
      code[1009] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010010011100001000000000000000000000000001000000011100011100000000001001101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1010] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100100110000000001000000101010000000000000000000000000000000000000000000100000000011010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1011] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1012] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010011100001000000000000000000000000000000000000000000100000000001001110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[1013] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010111110000000001011110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1014] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1015] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000010000000000000101110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1016] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1017] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000001010011100001000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[1018] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010101100000000001100000101010000000000000000000000000000000000000000000100000000101001110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1019] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011010011100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1020] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110011100001000000000000000000000000001000000010010101000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1021] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000001100110000000000000000101010000000000000000000000000001000000011010011000000000000000010101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[1022] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010110011100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1023] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001110011100001000000000000000000000000001000000010010101000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1024] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000011100110000000000000000101010000000000000000000000000001000000010110011000000000000000010101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[1025] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110011100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1026] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001011100001000000000000000000000000001000000000110101000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1027] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000000010110000000000000000101010000000000000000000000000001000000011110011100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[1028] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010001011100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1029] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001001011100001000000000000000000000000001000000000110101000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1030] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000010000000010010110000000000000000101010000000000000000000000000001000000010001011100000000001111001101000000000000000000000000000000000000000000010000000111011101000010000000000;                                          // moveLong
      code[1031] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1032] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100101010000000001000000101010000000000000000000000000000000000000000000100000000101011010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1033] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000001101010000000001000000101010000000000000000000000000000000000000000000100000000101011010000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1034] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001011100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1035] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000101011100001000000000000000000000000001000000011001011100000001110111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1036] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010101011100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1037] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001101011100001000000000000000000000000001000000010101011100000001110111001101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1038] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011101011100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1039] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000111010110000000000000000101010000000000000000000000000000000000000000000100000000010101110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1040] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000011011100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1041] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000000110110000000000000000101010000000000000000000000000000000000000000000100000000110101110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1042] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010011011100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1043] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000100110110000000000000000101010000000000000000000000000000000000000000000100000001001010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1044] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001011011100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1045] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010110110000000010000000101010000000000000000000000000000000000000000000100000000011010110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1046] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000010000000010101100000000000000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1047] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011011011100001000000000000000000000000001000000001010110000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1048] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000011011011100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000011000000000010000000000;                                          // resize
      code[1049] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000111011100001000000000000000000000000001000000001010110000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1050] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000000111011100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000111000000000010000000000;                                          // resize
      code[1051] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010111011100001000000000000000000000000001000000001010110000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1052] = 'b0000000000000000000000001000110000000000000000000000000000000000000000000000000000000000000000001000000010111011100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000100000000010000000000;                                          // resize
      code[1053] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000010000000000000011100110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1054] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000011000000000000010010110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1055] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1056] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001110100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1057] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000010010110100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1058] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1059] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011001110100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1060] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1061] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1062] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1063] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1064] = 'b0000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000001100000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // free
      code[1065] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000100100100000000001000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1066] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1067] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000101000100000000010111110100001000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000000010000000000010000000000;                                          // jNe
      code[1068] = 'b0000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000001000000001111011100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // in
      code[1069] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1070] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111011100001000000000000000000000000000000000011000000000000001100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1071] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000101000000000000001000001100001000000000000000000000000000000000000000000100000001111101110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jNe
      code[1072] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000100000001111101110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1073] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1074] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1075] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000111101000000000010000001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1076] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1077] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1078] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000000111100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1079] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1080] = 'b0000000000000000000000001001100000000000000000000000000000000000000000000000000000000000011001000000000001100001100001000000000000000000000000000000000000000000100000000000011110000100000000000000000000000000000000000000000000000000110001100000010000000000;                                          // jGe
      code[1081] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000001000000010000111100001000000000000000000000000001000000011111011000000000000000010101000000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[1082] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001000111100001000000000000000000000000001000000011111011000000000010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1083] = 'b0000000000000000000000001101100000000000000000000000000000000000000000000000000000000000101100000000000011100001100001000000000000000000000000000000000000000000100000000111101110000100000000000000000000000000100000000100011110000000100001110110100000000000;                                          // jLe
      code[1084] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011000111100001000000000000000000000000000000000000000000100000001000011110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[1085] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000001000000000100111100001000000000000000000000000001000000011111011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[1086] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000000010001100001000000000000000000000000000000000000000000100000000010011110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[1087] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000100000001111101110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1088] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1089] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000100000001100011110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1090] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000001000000000010000001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1091] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1092] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010100111100001000000000000000000000000001000000011111011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1093] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001100111100001000000000000000000000000001000000010100111100000001100011101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1094] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111011100001000000000000000000000000000000000000000000100000000110011110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1095] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001010000000000010100001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1096] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001110000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1097] = 'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000001000000011100111100001000000000000000000000000000000000000000000100000000100011110000100000000000000000000000000000000000000000010000000011110111000010000000000;                                          // arrayIndex
      code[1098] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000010010001100001000000000000000000000000000000000000000000100000001110011110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[1099] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000100000001111101110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1100] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1101] = 'b0000000000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000100000001110011110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // subtract
      code[1102] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001010000000000010000001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1103] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001001000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1104] = 'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000001000000000010111100001000000000000000000000000000000000000000000100000000100011110000100000000000000000000000000000000000000000010000000011110111000010000000000;                                          // arrayCountLess
      code[1105] = 'b0000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000001000000010010111100001000000000000000000000000001000000011111011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // not
      code[1106] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000001010001100001000000000000000000000000000000000000000000100000001001011110000100000000000000000000000000000000000000000000000000000000000000010000000000;                                          // jEq
      code[1107] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000100000001111101110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1108] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1109] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000100000000001011110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1110] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001100000000000010000001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1111] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1112] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001010111100001000000000000000000000000001000000011111011000000000110000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1113] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011010111100001000000000000000000000000001000000001010111100000000001011101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1114] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011111011100001000000000000000000000000000000000000000000100000001101011110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1115] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1116] = 'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000111100001000000000000000000000000000000000000000000100000000000011110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // add
      code[1117] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111111111010110110000000000100001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1118] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1119] = 'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // assert
      code[1120] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1121] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1122] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1123] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000110111100001000000000000000000000000000000000000000000000000001000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1124] = 'b0000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000100000000000011010001100001000000000000000000000000000000000000000000100000000011011110000100000000000000000000000000000000000000000000000000100000000000010000000000;                                          // jNe
      code[1125] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[1126] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000010110111100001000000000000000000000000000000000000000000000000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1127] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000001110111100001000000000000000000000000000000000000000000000000000100000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1128] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000011110111100001000000000000000000000000001000000010110111000000001010000010101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1129] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000001000000000001111100001000000000000000000000000001000000011110111100000000111011101101000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[1130] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000111110000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[1131] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000000110001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1132] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001101000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1133] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[1134] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000011000100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1135] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000001000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1136] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001011111000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1137] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000110000000000000011000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1138] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[1139] = 'b0000000000000000000000001111100000000000000000000000000000000000111111111111111111011111011100010000000010000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[1140] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
    end
  endtask

  task endTest();                                                               // BTree: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 0;
      success = success && outMem[1] == 1;
      success = success && outMem[2] == 22;
      success = success && outMem[3] == 0;
      success = success && outMem[4] == 1;
      success = success && outMem[5] == 33;
    end
  endtask
