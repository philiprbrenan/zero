//----------------------------------------------------------------------------
// NWayTree CPU
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2023
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module cpu(reset, next, clock, diA, doA, dI, dO, dcI, dcO, stop,                // The cpu executes one step in the computation per input clock. We can also put values into memory and get values out again to test each program.
  programCounter, rs, rt);
  input      reset;                                                             // Reset the cpu so that we can run the programs one after another
  input      next;                                                              // Run the next program
  input      clock;                                                             // Program counter
  input      dcI, dcO;                                                          // Data in and out clocks
  input [7:0]diA;                                                               // Data input address
  input [7:0]doA;                                                               // Data  output address
  input [7:0]dI;                                                                // Data input value
  output[7:0]dO;                                                                // Data output value
  output     stop;                                                              // Program has finished - stop was executed
  output [11:0]programCounter;                                                  // Program counter output
  output [15:0]rs;                                                              // Source register
  output [15:0]rt;                                                              // Target register
  always begin #1 $display("Memory in hex:"); end
  reg stopped;                                                                  // Set when we stop

//  reg [ 7:0] dia;                                                               // Data input address
  reg [ 7:0] doa;                                                               // Data output address

  reg [15:0] R [0:15];                                                          // Registers
  reg [ 7:0] D [0:2**8-1];                                                      // Data during program execution
  reg [ 7:0] DI[0:2**8-1];                                                      // Data as input - then copied to the actual data  at program start
  reg [ 7:0] DO[0:2**8-1];                                                      // Data as output - copied from actual memory after program execution
  reg [ 8:0] P [0:2**11-1];                                                     // Program

  reg [ 8:0] C;                                                                 // Constant
  reg [ 8:0] S;                                                                 // Source
  reg [ 8:0] T;                                                                 // Target

  integer pc = 0;                                                               // Program counter, next change in program counter
//  integer j = 0;                                                                // Jump target
  integer i = 0;                                                                // Current instruction
//  integer z = 0;                                                                // Instruction count
  integer idi, ido;                                                             // Input and output indices for data memeory
  integer iprogram = 0;                                                         // Number of the program to run

  integer resetN = 0, resetL = 0;
  integer nextN  = 0, nextL  = 0;

  assign dO   = DO[doa];                                                        // Assign the completed memory output value to the output pins
  assign stop = stopped > 0 ? 1 : 0;                                            // Show whether we have stopped yet or not
  assign programCounter = pc;                                                   // Show the program counter
  assign rs   = R[S];                                                           // Show the source register
  assign rt   = R[T];                                                           // Show the target register

  always @ (posedge dcI)   DI[diA]   <= dI;                                     // Write into data memory
  always @ (posedge dcO)   doa       <= doA;                                    // Read from data memory

  always @ (posedge reset) resetN <= resetN + 1;                                // Restart at the first program
  always @ (posedge next)  nextN   =  nextN + 1;                                // Run the next program

  always @ (posedge clock) begin                                                // Execute next step in program

    if (resetN != resetL) begin;                                                // Reset
      resetL <= resetN;
      iprogram <= 0;
      pc <= 0;
    end

    else if (nextN != nextL) begin;                                             // Next
      nextL <= nextN;

      R[0] = 0; R[1] = 0; R[ 2] = 0; R[ 3] = 0; R[ 4] = 0; R[ 5] = 0; R[ 6] = 0; R[ 7] = 0;
      R[8] = 0; R[9] = 0; R[10] = 0; R[11] = 0; R[12] = 0; R[13] = 0; R[14] = 0; R[15] = 0;

      for(idi = 0; idi < 2**8; idi = idi + 1) D[idi] = DI[idi];                // Load clocked in data

      C  <= 0;                                                                  // Clear constant box
      S  <= 0;                                                                  // Clear source box
      T  <= 0;                                                                  // Clear target box

      if (iprogram == 0) load_Program1;                                         // Load program 1
      if (iprogram == 1) load_Program2;                                         // Load program 2
      if (iprogram == 2) load_Program3;                                         // Load program 3
      if (iprogram == 3) load_Instructions;                                     // Load test programs
      if (iprogram == 4) load_1_to_3;
      if (iprogram == 5) load_For_Loop;
      if (iprogram == 6) load_If;
      if (iprogram == 7) load_ParityBits;

      iprogram <= iprogram + 1;                                                 // Select the next program

      stopped <= 0;                                                             // We are now executing the program so we are not stopped
      pc <= 0;                                                                  // Start at the first instruction allowing for the clock going negative
    end

    else if (P[pc] <= 9'b0_1111_1111) begin; C <= P[pc];                  ppc(); end  // Constant
    else if (P[pc] <= 9'b1_0111_1111) begin; S <= P[pc] & 9'b0_0011_1111; ppc(); end  // Source
    else if (P[pc] <= 9'b1_1011_1111) begin; T <= P[pc] & 9'b0_0011_1111; ppc(); end  // Target
    else begin                                                                        // Decode opcode
      case(P[pc] & 6'h1f)
         0 : begin; R[T]    <=   rt  + rs;                                ppc(); end  // add
         1 : begin; R[T]    <=   rt  & rs;                                ppc(); end  // and
         2 : begin; R[T]    <=   rs == rt ? 1 : 0;                        ppc(); end  // cmpEq
         3 : begin; R[S]    <=   rs  >   C  ? 1 : 0;                      ppc(); end  // cmpGt
         4 : begin; R[S]    <=   rs  <   C  ? 1 : 0;                      ppc(); end  // cmpLt
         5 : begin; R[S]    <=   rs  - 1;                                 ppc(); end  // dec
         6 : begin; R[S]    <=   rs  + 1;                                 ppc(); end  // inc
         7 : begin; pc      <=   rs  > 0    ? (C << 3 ) - 2 : pc + 1;            end  // jumpIfNotZero - the minus three compensates for the fact that we are going to increment the program counter
         8 : begin; pc      <=   rs == 0    ? (C << 3 ) - 2 : pc + 1;            end  // jumpIfZero
         9 : begin; ppc();                                                       end  // label
        10 : begin; R[S]    <=   C;                                       ppc(); end  // ldrc
        11 : begin; R[S]    <=   D[C];                                    ppc(); end  // ldrd
        12 : begin; R[T]    <=   D[rs];                                   ppc(); end  // ldri
        13 : begin; R[T]    <=   rs;                                      ppc(); end  // ldrr
        14 : begin; R[S]    <= ! rs;                                      ppc(); end  // not
        15 : begin; R[T]    <=   rt | rs;                                 ppc(); end  // or
        16 : begin; R[S]    <=   rs << C;                                 ppc(); end  // sl
        17 : begin; R[S]    <=   rs >> C;                                 ppc(); end  // sr
        18 : begin; D[C]    <=   rs;                                      ppc(); end  // strd
        19 : begin; D[R[S]] <=   rt;                                      ppc(); end  // stri
        20 : begin; R[T]    <=   rt  - rs;                                ppc(); end  // sub
        21 : begin; R[S]    <=   rs  ^   C;                               ppc(); end  // xor
        22 : begin                                                                   // stop
          //$display("Memory in decimal:");
          //for(i = 0; i < 2**8; i = i + 16) begin                                // Print memory in decimal
          //  $display(i, " ", D[i+0], " ", D[i+1], " ", D[i+2], " ", D[i+3], "  ", D[i+4], " ", D[i+5], " ", D[i+6], " ", D[i+7], "   ", D[i+8], " ", D[i+9], " ", D[i+10], " ", D[i+11], "  ", D[i+12], " ", D[i+13], " ", D[i+14], " ", D[i+15]);
          //end
          //$display("Memory in hex:");
          //for(i = 0; i < 2**8; i = i + 16) begin                                // Print memory in hexadecimal
          //  $displayh(i, " ", D[i+0], " ", D[i+1], " ", D[i+2], " ", D[i+3], "  ", D[i+4], " ", D[i+5], " ", D[i+6], " ", D[i+7], "   ", D[i+8], " ", D[i+9], " ", D[i+10], " ", D[i+11], "  ", D[i+12], " ", D[i+13], " ", D[i+14], " ", D[i+15]);
          //end
          //$display("Finished");
          for(ido = 0; ido < 2**8; ido = ido + 1) DO[ido] <= D[ido];            // Place data in output area
          stopped <= 1;
        end
      endcase
    end
  end

  task ppc;                                                                     // Increment program counter
    begin
      pc <= pc + 1;
    end
  endtask

//  always @ (negedge clock) begin                                              // Trace program execution
//    $displayh("%08d  %05d   %8x   %3x %3x %3x   %4x %4x %4x %4x   %4x %4x %4x %4x     %4x %4x %4x %4x   %4x %4x %4x %4x",
//        z, pc, i,   C, S, T, R[0], R[1], R[2], R[3], R[4], R[5], R[6], R[7], R[8], R[9], R[10], R[11], R[12], R[13], R[14], R[15]);
//    z = z + 1;
//  end

  task  automatic load_Instructions;                                                       // Load instructions
    begin
      $display("Instructions");
      P[   0] <= 9'b000000001; // Load the constant box with 1
      P[   1] <= 9'b101001110; // Load the source box with 14
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   4] <= 9'b000000010; // Load the constant box with 2
      P[   5] <= 9'b101001111; // Load the source box with 15
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   8] <= 9'b000000000; // Load the constant box with 0
      P[   9] <= 9'b101001111; // Load the source box with 15
      P[  10] <= 9'b110001110; // Load the target box with 14
      P[  11] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[  12] <= 9'b000000000; // Load the constant box with 0
      P[  13] <= 9'b101001110; // Load the source box with 14
      P[  14] <= 9'b110000000; // Load the target box with 0
      P[  15] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  16] <= 9'b000010101; // Load the constant box with 21
      P[  17] <= 9'b101001111; // Load the source box with 15
      P[  18] <= 9'b110000000; // Load the target box with 0
      P[  19] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  20] <= 9'b000000000; // Load the constant box with 0
      P[  21] <= 9'b101001111; // Load the source box with 15
      P[  22] <= 9'b110000000; // Load the target box with 0
      P[  23] <= 9'b111001110; // not: Invert the bits in a register
      P[  24] <= 9'b000000001; // Load the constant box with 1
      P[  25] <= 9'b101001111; // Load the source box with 15
      P[  26] <= 9'b110000000; // Load the target box with 0
      P[  27] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  28] <= 9'b000000101; // Load the constant box with 5
      P[  29] <= 9'b101001110; // Load the source box with 14
      P[  30] <= 9'b110000000; // Load the target box with 0
      P[  31] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  32] <= 9'b000001001; // Load the constant box with 9
      P[  33] <= 9'b101001111; // Load the source box with 15
      P[  34] <= 9'b110000000; // Load the target box with 0
      P[  35] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  36] <= 9'b000000000; // Load the constant box with 0
      P[  37] <= 9'b101001111; // Load the source box with 15
      P[  38] <= 9'b110001110; // Load the target box with 14
      P[  39] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[  40] <= 9'b000000010; // Load the constant box with 2
      P[  41] <= 9'b101001110; // Load the source box with 14
      P[  42] <= 9'b110000000; // Load the target box with 0
      P[  43] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  44] <= 9'b000000101; // Load the constant box with 5
      P[  45] <= 9'b101001110; // Load the source box with 14
      P[  46] <= 9'b110000000; // Load the target box with 0
      P[  47] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  48] <= 9'b000001001; // Load the constant box with 9
      P[  49] <= 9'b101001111; // Load the source box with 15
      P[  50] <= 9'b110000000; // Load the target box with 0
      P[  51] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  52] <= 9'b000000000; // Load the constant box with 0
      P[  53] <= 9'b101001111; // Load the source box with 15
      P[  54] <= 9'b110001110; // Load the target box with 14
      P[  55] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[  56] <= 9'b000000011; // Load the constant box with 3
      P[  57] <= 9'b101001110; // Load the source box with 14
      P[  58] <= 9'b110000000; // Load the target box with 0
      P[  59] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  60] <= 9'b000010101; // Load the constant box with 21
      P[  61] <= 9'b101000010; // Load the source box with 2
      P[  62] <= 9'b110000000; // Load the target box with 0
      P[  63] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  64] <= 9'b000000000; // Load the constant box with 0
      P[  65] <= 9'b101000010; // Load the source box with 2
      P[  66] <= 9'b110000000; // Load the target box with 0
      P[  67] <= 9'b111000110; // inc: Increment a register by one
      P[  68] <= 9'b000000100; // Load the constant box with 4
      P[  69] <= 9'b101000010; // Load the source box with 2
      P[  70] <= 9'b110000000; // Load the target box with 0
      P[  71] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  72] <= 9'b000000000; // Load the constant box with 0
      P[  73] <= 9'b101000010; // Load the source box with 2
      P[  74] <= 9'b110000011; // Load the target box with 3
      P[  75] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  76] <= 9'b000000000; // Load the constant box with 0
      P[  77] <= 9'b101000011; // Load the source box with 3
      P[  78] <= 9'b110000000; // Load the target box with 0
      P[  79] <= 9'b111000101; // dec: Decrement a register by one
      P[  80] <= 9'b000000101; // Load the constant box with 5
      P[  81] <= 9'b101000011; // Load the source box with 3
      P[  82] <= 9'b110000000; // Load the target box with 0
      P[  83] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  84] <= 9'b000000011; // Load the constant box with 3
      P[  85] <= 9'b101000010; // Load the source box with 2
      P[  86] <= 9'b110000000; // Load the target box with 0
      P[  87] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  88] <= 9'b000000001; // Load the constant box with 1
      P[  89] <= 9'b101000010; // Load the source box with 2
      P[  90] <= 9'b110000000; // Load the target box with 0
      P[  91] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  92] <= 9'b000000110; // Load the constant box with 6
      P[  93] <= 9'b101000010; // Load the source box with 2
      P[  94] <= 9'b110000000; // Load the target box with 0
      P[  95] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  96] <= 9'b000000011; // Load the constant box with 3
      P[  97] <= 9'b101000010; // Load the source box with 2
      P[  98] <= 9'b110000000; // Load the target box with 0
      P[  99] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 100] <= 9'b000000010; // Load the constant box with 2
      P[ 101] <= 9'b101000010; // Load the source box with 2
      P[ 102] <= 9'b110000000; // Load the target box with 0
      P[ 103] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 104] <= 9'b000000111; // Load the constant box with 7
      P[ 105] <= 9'b101000010; // Load the source box with 2
      P[ 106] <= 9'b110000000; // Load the target box with 0
      P[ 107] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 108] <= 9'b000010100; // Load the constant box with 20
      P[ 109] <= 9'b101000100; // Load the source box with 4
      P[ 110] <= 9'b110000000; // Load the target box with 0
      P[ 111] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 112] <= 9'b000001001; // Load the constant box with 9
      P[ 113] <= 9'b101000101; // Load the source box with 5
      P[ 114] <= 9'b110000000; // Load the target box with 0
      P[ 115] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 116] <= 9'b000000000; // Load the constant box with 0
      P[ 117] <= 9'b101000101; // Load the source box with 5
      P[ 118] <= 9'b110000100; // Load the target box with 4
      P[ 119] <= 9'b111010100; // sub: Subtract the second register from the first register replace the first register with the result
      P[ 120] <= 9'b000001000; // Load the constant box with 8
      P[ 121] <= 9'b101000100; // Load the source box with 4
      P[ 122] <= 9'b110000000; // Load the target box with 0
      P[ 123] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 124] <= 9'b000001001; // Load the constant box with 9
      P[ 125] <= 9'b101000001; // Load the source box with 1
      P[ 126] <= 9'b110000000; // Load the target box with 0
      P[ 127] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 128] <= 9'b001100011; // Load the constant box with 99
      P[ 129] <= 9'b101000010; // Load the source box with 2
      P[ 130] <= 9'b110000000; // Load the target box with 0
      P[ 131] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 132] <= 9'b000000000; // Load the constant box with 0
      P[ 133] <= 9'b101000001; // Load the source box with 1
      P[ 134] <= 9'b110000010; // Load the target box with 2
      P[ 135] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[ 136] <= 9'b000000000; // Load the constant box with 0
      P[ 137] <= 9'b101000000; // Load the source box with 0
      P[ 138] <= 9'b110000000; // Load the target box with 0
      P[ 139] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task  automatic load_1_to_3;                                                             // Test program
    begin
      $display("Program 1_to_3");
      P[     0] <= 9'b000000000; // Load the constant box with 0
      P[     1] <= 9'b101000000; // Load the source box with 0
      P[     2] <= 9'b110000000; // Load the target box with 0
      P[     3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[     4] <= 9'b000000000; // Load the constant box with 0
      P[     5] <= 9'b101000000; // Load the source box with 0
      P[     6] <= 9'b110000000; // Load the target box with 0
      P[     7] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[     8] <= 9'b000000000; // Load the constant box with 0
      P[     9] <= 9'b101000000; // Load the source box with 0
      P[    10] <= 9'b110000000; // Load the target box with 0
      P[    11] <= 9'b111000110; // inc: Increment a register by one
      P[    12] <= 9'b000000001; // Load the constant box with 1
      P[    13] <= 9'b101000000; // Load the source box with 0
      P[    14] <= 9'b110000000; // Load the target box with 0
      P[    15] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[    16] <= 9'b000000000; // Load the constant box with 0
      P[    17] <= 9'b101000000; // Load the source box with 0
      P[    18] <= 9'b110000000; // Load the target box with 0
      P[    19] <= 9'b111000110; // inc: Increment a register by one
      P[    20] <= 9'b000000010; // Load the constant box with 2
      P[    21] <= 9'b101000000; // Load the source box with 0
      P[    22] <= 9'b110000000; // Load the target box with 0
      P[    23] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[    24] <= 9'b000000000; // Load the constant box with 0
      P[    25] <= 9'b101000000; // Load the source box with 0
      P[    26] <= 9'b110000000; // Load the target box with 0
      P[    27] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task  automatic load_For_Loop;                                                           // For Loop low
    begin
      $display("Program For_Loop");
      P[   0] <= 9'b011111111; // Load the constant box with 255
      P[   1] <= 9'b101000000; // Load the source box with 0
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   4] <= 9'b000000001; // Load the constant box with 1
      P[   5] <= 9'b101000000; // Load the source box with 0
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001001; // label: Create and set a label
      P[   8] <= 9'b000000000; // Load the constant box with 0
      P[   9] <= 9'b101000000; // Load the source box with 0
      P[  10] <= 9'b110000000; // Load the target box with 0
      P[  11] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[  12] <= 9'b000000000; // Load the constant box with 0
      P[  13] <= 9'b101000000; // Load the source box with 0
      P[  14] <= 9'b110000000; // Load the target box with 0
      P[  15] <= 9'b111000101; // dec: Decrement a register by one
      P[  16] <= 9'b000000001; // Load the constant box with 1
      P[  17] <= 9'b101000000; // Load the source box with 0
      P[  18] <= 9'b110000000; // Load the target box with 0
      P[  19] <= 9'b111000111; // jumpIfNotZero: Jump backwards to the specified location in the program if the register is not zero - useful for constructing for loops
      P[  20] <= 9'b000000000; // Load the constant box with 0
      P[  21] <= 9'b101000000; // Load the source box with 0
      P[  22] <= 9'b110000000; // Load the target box with 0
      P[  23] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task  automatic load_If;                                                                 // If low
    begin
      $display("Program If");
      P[   0] <= 9'b011111111; // Load the constant box with 255
      P[   1] <= 9'b101000000; // Load the source box with 0
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   4] <= 9'b000000010; // Load the constant box with 2
      P[   5] <= 9'b101000000; // Load the source box with 0
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001001; // label: Create and set a label
      P[   8] <= 9'b000000000; // Load the constant box with 0
      P[   9] <= 9'b101000000; // Load the source box with 0
      P[  10] <= 9'b110000001; // Load the target box with 1
      P[  11] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  12] <= 9'b000001111; // Load the constant box with 15
      P[  13] <= 9'b101000001; // Load the source box with 1
      P[  14] <= 9'b110000000; // Load the target box with 0
      P[  15] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  16] <= 9'b000001111; // Load the constant box with 15
      P[  17] <= 9'b101000001; // Load the source box with 1
      P[  18] <= 9'b110000000; // Load the target box with 0
      P[  19] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  20] <= 9'b000000100; // Load the constant box with 4
      P[  21] <= 9'b101000001; // Load the source box with 1
      P[  22] <= 9'b110000000; // Load the target box with 0
      P[  23] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[  24] <= 9'b000000000; // Load the constant box with 0
      P[  25] <= 9'b101000000; // Load the source box with 0
      P[  26] <= 9'b110000000; // Load the target box with 0
      P[  27] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[  28] <= 9'b000000010; // Load the constant box with 2
      P[  29] <= 9'b101000000; // Load the source box with 0
      P[  30] <= 9'b110000000; // Load the target box with 0
      P[  31] <= 9'b111001001; // label: Set a label
      P[  32] <= 9'b000000000; // Load the constant box with 0
      P[  33] <= 9'b101000000; // Load the source box with 0
      P[  34] <= 9'b110000000; // Load the target box with 0
      P[  35] <= 9'b111000101; // dec: Decrement a register by one
      P[  36] <= 9'b000000001; // Load the constant box with 1
      P[  37] <= 9'b101000000; // Load the source box with 0
      P[  38] <= 9'b110000000; // Load the target box with 0
      P[  39] <= 9'b111000111; // jumpIfNotZero: Jump backwards to the specified location in the program if the register is not zero - useful for constructing for loops
      P[  40] <= 9'b000000000; // Load the constant box with 0
      P[  41] <= 9'b101000000; // Load the source box with 0
      P[  42] <= 9'b110000000; // Load the target box with 0
      P[  43] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task automatic load_ParityBits;                                                         // ParityBits
    begin
      $display("ParityBits");
      P[   0] <= 9'b011111110; // Load the constant box with 254
      P[   1] <= 9'b101000001; // Load the source box with 1
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[   4] <= 9'b011111101; // Load the constant box with 253
      P[   5] <= 9'b101000010; // Load the source box with 2
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[   8] <= 9'b000001000; // Load the constant box with 8
      P[   9] <= 9'b101000001; // Load the source box with 1
      P[  10] <= 9'b110000000; // Load the target box with 0
      P[  11] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  12] <= 9'b000000000; // Load the constant box with 0
      P[  13] <= 9'b101000010; // Load the source box with 2
      P[  14] <= 9'b110000001; // Load the target box with 1
      P[  15] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[  16] <= 9'b000000000; // Load the constant box with 0
      P[  17] <= 9'b101000001; // Load the source box with 1
      P[  18] <= 9'b110000010; // Load the target box with 2
      P[  19] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  20] <= 9'b000000101; // Load the constant box with 5
      P[  21] <= 9'b101000010; // Load the source box with 2
      P[  22] <= 9'b110000000; // Load the target box with 0
      P[  23] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  24] <= 9'b000001111; // Load the constant box with 15
      P[  25] <= 9'b101000010; // Load the source box with 2
      P[  26] <= 9'b110000000; // Load the target box with 0
      P[  27] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  28] <= 9'b000000000; // Load the constant box with 0
      P[  29] <= 9'b101000001; // Load the source box with 1
      P[  30] <= 9'b110000011; // Load the target box with 3
      P[  31] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  32] <= 9'b000000110; // Load the constant box with 6
      P[  33] <= 9'b101000011; // Load the source box with 3
      P[  34] <= 9'b110000000; // Load the target box with 0
      P[  35] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  36] <= 9'b000001111; // Load the constant box with 15
      P[  37] <= 9'b101000011; // Load the source box with 3
      P[  38] <= 9'b110000000; // Load the target box with 0
      P[  39] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  40] <= 9'b000000000; // Load the constant box with 0
      P[  41] <= 9'b101000001; // Load the source box with 1
      P[  42] <= 9'b110000100; // Load the target box with 4
      P[  43] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  44] <= 9'b000000111; // Load the constant box with 7
      P[  45] <= 9'b101000100; // Load the source box with 4
      P[  46] <= 9'b110000000; // Load the target box with 0
      P[  47] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  48] <= 9'b000001111; // Load the constant box with 15
      P[  49] <= 9'b101000100; // Load the source box with 4
      P[  50] <= 9'b110000000; // Load the target box with 0
      P[  51] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  52] <= 9'b000000000; // Load the constant box with 0
      P[  53] <= 9'b101000001; // Load the source box with 1
      P[  54] <= 9'b110000101; // Load the target box with 5
      P[  55] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  56] <= 9'b000001000; // Load the constant box with 8
      P[  57] <= 9'b101000101; // Load the source box with 5
      P[  58] <= 9'b110000000; // Load the target box with 0
      P[  59] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  60] <= 9'b000001111; // Load the constant box with 15
      P[  61] <= 9'b101000101; // Load the source box with 5
      P[  62] <= 9'b110000000; // Load the target box with 0
      P[  63] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  64] <= 9'b000000000; // Load the constant box with 0
      P[  65] <= 9'b101000001; // Load the source box with 1
      P[  66] <= 9'b110000110; // Load the target box with 6
      P[  67] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  68] <= 9'b000001001; // Load the constant box with 9
      P[  69] <= 9'b101000110; // Load the source box with 6
      P[  70] <= 9'b110000000; // Load the target box with 0
      P[  71] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  72] <= 9'b000001111; // Load the constant box with 15
      P[  73] <= 9'b101000110; // Load the source box with 6
      P[  74] <= 9'b110000000; // Load the target box with 0
      P[  75] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  76] <= 9'b000000000; // Load the constant box with 0
      P[  77] <= 9'b101000001; // Load the source box with 1
      P[  78] <= 9'b110000111; // Load the target box with 7
      P[  79] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  80] <= 9'b000001010; // Load the constant box with 10
      P[  81] <= 9'b101000111; // Load the source box with 7
      P[  82] <= 9'b110000000; // Load the target box with 0
      P[  83] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  84] <= 9'b000001111; // Load the constant box with 15
      P[  85] <= 9'b101000111; // Load the source box with 7
      P[  86] <= 9'b110000000; // Load the target box with 0
      P[  87] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  88] <= 9'b000000000; // Load the constant box with 0
      P[  89] <= 9'b101000001; // Load the source box with 1
      P[  90] <= 9'b110001000; // Load the target box with 8
      P[  91] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  92] <= 9'b000001011; // Load the constant box with 11
      P[  93] <= 9'b101001000; // Load the source box with 8
      P[  94] <= 9'b110000000; // Load the target box with 0
      P[  95] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  96] <= 9'b000001111; // Load the constant box with 15
      P[  97] <= 9'b101001000; // Load the source box with 8
      P[  98] <= 9'b110000000; // Load the target box with 0
      P[  99] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 100] <= 9'b000000000; // Load the constant box with 0
      P[ 101] <= 9'b101000001; // Load the source box with 1
      P[ 102] <= 9'b110001001; // Load the target box with 9
      P[ 103] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 104] <= 9'b000001100; // Load the constant box with 12
      P[ 105] <= 9'b101001001; // Load the source box with 9
      P[ 106] <= 9'b110000000; // Load the target box with 0
      P[ 107] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 108] <= 9'b000001111; // Load the constant box with 15
      P[ 109] <= 9'b101001001; // Load the source box with 9
      P[ 110] <= 9'b110000000; // Load the target box with 0
      P[ 111] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 112] <= 9'b000000000; // Load the constant box with 0
      P[ 113] <= 9'b101000001; // Load the source box with 1
      P[ 114] <= 9'b110001010; // Load the target box with 10
      P[ 115] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 116] <= 9'b000001101; // Load the constant box with 13
      P[ 117] <= 9'b101001010; // Load the source box with 10
      P[ 118] <= 9'b110000000; // Load the target box with 0
      P[ 119] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 120] <= 9'b000001111; // Load the constant box with 15
      P[ 121] <= 9'b101001010; // Load the source box with 10
      P[ 122] <= 9'b110000000; // Load the target box with 0
      P[ 123] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 124] <= 9'b000000000; // Load the constant box with 0
      P[ 125] <= 9'b101000001; // Load the source box with 1
      P[ 126] <= 9'b110001011; // Load the target box with 11
      P[ 127] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 128] <= 9'b000001110; // Load the constant box with 14
      P[ 129] <= 9'b101001011; // Load the source box with 11
      P[ 130] <= 9'b110000000; // Load the target box with 0
      P[ 131] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 132] <= 9'b000001111; // Load the constant box with 15
      P[ 133] <= 9'b101001011; // Load the source box with 11
      P[ 134] <= 9'b110000000; // Load the target box with 0
      P[ 135] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 136] <= 9'b000000000; // Load the constant box with 0
      P[ 137] <= 9'b101000001; // Load the source box with 1
      P[ 138] <= 9'b110001100; // Load the target box with 12
      P[ 139] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 140] <= 9'b000001111; // Load the constant box with 15
      P[ 141] <= 9'b101001100; // Load the source box with 12
      P[ 142] <= 9'b110000000; // Load the target box with 0
      P[ 143] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 144] <= 9'b000001111; // Load the constant box with 15
      P[ 145] <= 9'b101001100; // Load the source box with 12
      P[ 146] <= 9'b110000000; // Load the target box with 0
      P[ 147] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 148] <= 9'b000000000; // Load the constant box with 0
      P[ 149] <= 9'b101000001; // Load the source box with 1
      P[ 150] <= 9'b110001101; // Load the target box with 13
      P[ 151] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 152] <= 9'b000000101; // Load the constant box with 5
      P[ 153] <= 9'b101001101; // Load the source box with 13
      P[ 154] <= 9'b110000000; // Load the target box with 0
      P[ 155] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 156] <= 9'b000001001; // Load the constant box with 9
      P[ 157] <= 9'b101001101; // Load the source box with 13
      P[ 158] <= 9'b110000000; // Load the target box with 0
      P[ 159] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 160] <= 9'b000000001; // Load the constant box with 1
      P[ 161] <= 9'b101001101; // Load the source box with 13
      P[ 162] <= 9'b110000000; // Load the target box with 0
      P[ 163] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 164] <= 9'b000000000; // Load the constant box with 0
      P[ 165] <= 9'b101000001; // Load the source box with 1
      P[ 166] <= 9'b110001110; // Load the target box with 14
      P[ 167] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 168] <= 9'b000001000; // Load the constant box with 8
      P[ 169] <= 9'b101001110; // Load the source box with 14
      P[ 170] <= 9'b110000000; // Load the target box with 0
      P[ 171] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 172] <= 9'b000001101; // Load the constant box with 13
      P[ 173] <= 9'b101001110; // Load the source box with 14
      P[ 174] <= 9'b110000000; // Load the target box with 0
      P[ 175] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 176] <= 9'b000000101; // Load the constant box with 5
      P[ 177] <= 9'b101001110; // Load the source box with 14
      P[ 178] <= 9'b110000000; // Load the target box with 0
      P[ 179] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 180] <= 9'b000000000; // Load the constant box with 0
      P[ 181] <= 9'b101000001; // Load the source box with 1
      P[ 182] <= 9'b110001111; // Load the target box with 15
      P[ 183] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 184] <= 9'b000001111; // Load the constant box with 15
      P[ 185] <= 9'b101001111; // Load the source box with 15
      P[ 186] <= 9'b110000000; // Load the target box with 0
      P[ 187] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 188] <= 9'b000001100; // Load the constant box with 12
      P[ 189] <= 9'b101001111; // Load the source box with 15
      P[ 190] <= 9'b110000000; // Load the target box with 0
      P[ 191] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 192] <= 9'b000000000; // Load the constant box with 0
      P[ 193] <= 9'b101001111; // Load the source box with 15
      P[ 194] <= 9'b110001110; // Load the target box with 14
      P[ 195] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 196] <= 9'b000000000; // Load the constant box with 0
      P[ 197] <= 9'b101000010; // Load the source box with 2
      P[ 198] <= 9'b110001111; // Load the target box with 15
      P[ 199] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 200] <= 9'b000000000; // Load the constant box with 0
      P[ 201] <= 9'b101000011; // Load the source box with 3
      P[ 202] <= 9'b110001111; // Load the target box with 15
      P[ 203] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 204] <= 9'b000000000; // Load the constant box with 0
      P[ 205] <= 9'b101000100; // Load the source box with 4
      P[ 206] <= 9'b110001111; // Load the target box with 15
      P[ 207] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 208] <= 9'b000000000; // Load the constant box with 0
      P[ 209] <= 9'b101000101; // Load the source box with 5
      P[ 210] <= 9'b110001111; // Load the target box with 15
      P[ 211] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 212] <= 9'b000000000; // Load the constant box with 0
      P[ 213] <= 9'b101000110; // Load the source box with 6
      P[ 214] <= 9'b110001111; // Load the target box with 15
      P[ 215] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 216] <= 9'b000000000; // Load the constant box with 0
      P[ 217] <= 9'b101000111; // Load the source box with 7
      P[ 218] <= 9'b110001111; // Load the target box with 15
      P[ 219] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 220] <= 9'b000000000; // Load the constant box with 0
      P[ 221] <= 9'b101001000; // Load the source box with 8
      P[ 222] <= 9'b110001111; // Load the target box with 15
      P[ 223] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 224] <= 9'b000000001; // Load the constant box with 1
      P[ 225] <= 9'b101000000; // Load the source box with 0
      P[ 226] <= 9'b110000000; // Load the target box with 0
      P[ 227] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 228] <= 9'b000000000; // Load the constant box with 0
      P[ 229] <= 9'b101001111; // Load the source box with 15
      P[ 230] <= 9'b110000000; // Load the target box with 0
      P[ 231] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 232] <= 9'b011110111; // Load the constant box with 247
      P[ 233] <= 9'b101000000; // Load the source box with 0
      P[ 234] <= 9'b110000000; // Load the target box with 0
      P[ 235] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 236] <= 9'b000000000; // Load the constant box with 0
      P[ 237] <= 9'b101000000; // Load the source box with 0
      P[ 238] <= 9'b110000001; // Load the target box with 1
      P[ 239] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 240] <= 9'b000000000; // Load the constant box with 0
      P[ 241] <= 9'b101000000; // Load the source box with 0
      P[ 242] <= 9'b110001101; // Load the target box with 13
      P[ 243] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 244] <= 9'b000000000; // Load the constant box with 0
      P[ 245] <= 9'b101000010; // Load the source box with 2
      P[ 246] <= 9'b110001111; // Load the target box with 15
      P[ 247] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 248] <= 9'b000000000; // Load the constant box with 0
      P[ 249] <= 9'b101000011; // Load the source box with 3
      P[ 250] <= 9'b110001111; // Load the target box with 15
      P[ 251] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 252] <= 9'b000000000; // Load the constant box with 0
      P[ 253] <= 9'b101000100; // Load the source box with 4
      P[ 254] <= 9'b110001111; // Load the target box with 15
      P[ 255] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 256] <= 9'b000000000; // Load the constant box with 0
      P[ 257] <= 9'b101000101; // Load the source box with 5
      P[ 258] <= 9'b110001111; // Load the target box with 15
      P[ 259] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 260] <= 9'b000000000; // Load the constant box with 0
      P[ 261] <= 9'b101001001; // Load the source box with 9
      P[ 262] <= 9'b110001111; // Load the target box with 15
      P[ 263] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 264] <= 9'b000000000; // Load the constant box with 0
      P[ 265] <= 9'b101001010; // Load the source box with 10
      P[ 266] <= 9'b110001111; // Load the target box with 15
      P[ 267] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 268] <= 9'b000000000; // Load the constant box with 0
      P[ 269] <= 9'b101001011; // Load the source box with 11
      P[ 270] <= 9'b110001111; // Load the target box with 15
      P[ 271] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 272] <= 9'b000000001; // Load the constant box with 1
      P[ 273] <= 9'b101000000; // Load the source box with 0
      P[ 274] <= 9'b110000000; // Load the target box with 0
      P[ 275] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 276] <= 9'b000000000; // Load the constant box with 0
      P[ 277] <= 9'b101001111; // Load the source box with 15
      P[ 278] <= 9'b110000000; // Load the target box with 0
      P[ 279] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 280] <= 9'b011111000; // Load the constant box with 248
      P[ 281] <= 9'b101000000; // Load the source box with 0
      P[ 282] <= 9'b110000000; // Load the target box with 0
      P[ 283] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 284] <= 9'b000000000; // Load the constant box with 0
      P[ 285] <= 9'b101000000; // Load the source box with 0
      P[ 286] <= 9'b110000001; // Load the target box with 1
      P[ 287] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 288] <= 9'b000000100; // Load the constant box with 4
      P[ 289] <= 9'b101000000; // Load the source box with 0
      P[ 290] <= 9'b110000000; // Load the target box with 0
      P[ 291] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 292] <= 9'b000000000; // Load the constant box with 0
      P[ 293] <= 9'b101000000; // Load the source box with 0
      P[ 294] <= 9'b110001110; // Load the target box with 14
      P[ 295] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 296] <= 9'b000000000; // Load the constant box with 0
      P[ 297] <= 9'b101000010; // Load the source box with 2
      P[ 298] <= 9'b110001111; // Load the target box with 15
      P[ 299] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 300] <= 9'b000000000; // Load the constant box with 0
      P[ 301] <= 9'b101000011; // Load the source box with 3
      P[ 302] <= 9'b110001111; // Load the target box with 15
      P[ 303] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 304] <= 9'b000000000; // Load the constant box with 0
      P[ 305] <= 9'b101000110; // Load the source box with 6
      P[ 306] <= 9'b110001111; // Load the target box with 15
      P[ 307] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 308] <= 9'b000000000; // Load the constant box with 0
      P[ 309] <= 9'b101000111; // Load the source box with 7
      P[ 310] <= 9'b110001111; // Load the target box with 15
      P[ 311] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 312] <= 9'b000000000; // Load the constant box with 0
      P[ 313] <= 9'b101001001; // Load the source box with 9
      P[ 314] <= 9'b110001111; // Load the target box with 15
      P[ 315] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 316] <= 9'b000000000; // Load the constant box with 0
      P[ 317] <= 9'b101001010; // Load the source box with 10
      P[ 318] <= 9'b110001111; // Load the target box with 15
      P[ 319] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 320] <= 9'b000000000; // Load the constant box with 0
      P[ 321] <= 9'b101001100; // Load the source box with 12
      P[ 322] <= 9'b110001111; // Load the target box with 15
      P[ 323] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 324] <= 9'b000000001; // Load the constant box with 1
      P[ 325] <= 9'b101000000; // Load the source box with 0
      P[ 326] <= 9'b110000000; // Load the target box with 0
      P[ 327] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 328] <= 9'b000000000; // Load the constant box with 0
      P[ 329] <= 9'b101001111; // Load the source box with 15
      P[ 330] <= 9'b110000000; // Load the target box with 0
      P[ 331] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 332] <= 9'b011111001; // Load the constant box with 249
      P[ 333] <= 9'b101000000; // Load the source box with 0
      P[ 334] <= 9'b110000000; // Load the target box with 0
      P[ 335] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 336] <= 9'b000000000; // Load the constant box with 0
      P[ 337] <= 9'b101000000; // Load the source box with 0
      P[ 338] <= 9'b110000001; // Load the target box with 1
      P[ 339] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 340] <= 9'b000000010; // Load the constant box with 2
      P[ 341] <= 9'b101000000; // Load the source box with 0
      P[ 342] <= 9'b110000000; // Load the target box with 0
      P[ 343] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 344] <= 9'b000000000; // Load the constant box with 0
      P[ 345] <= 9'b101000000; // Load the source box with 0
      P[ 346] <= 9'b110001110; // Load the target box with 14
      P[ 347] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 348] <= 9'b000000000; // Load the constant box with 0
      P[ 349] <= 9'b101000010; // Load the source box with 2
      P[ 350] <= 9'b110001111; // Load the target box with 15
      P[ 351] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 352] <= 9'b000000000; // Load the constant box with 0
      P[ 353] <= 9'b101000100; // Load the source box with 4
      P[ 354] <= 9'b110001111; // Load the target box with 15
      P[ 355] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 356] <= 9'b000000000; // Load the constant box with 0
      P[ 357] <= 9'b101000110; // Load the source box with 6
      P[ 358] <= 9'b110001111; // Load the target box with 15
      P[ 359] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 360] <= 9'b000000000; // Load the constant box with 0
      P[ 361] <= 9'b101001000; // Load the source box with 8
      P[ 362] <= 9'b110001111; // Load the target box with 15
      P[ 363] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 364] <= 9'b000000000; // Load the constant box with 0
      P[ 365] <= 9'b101001001; // Load the source box with 9
      P[ 366] <= 9'b110001111; // Load the target box with 15
      P[ 367] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 368] <= 9'b000000000; // Load the constant box with 0
      P[ 369] <= 9'b101001011; // Load the source box with 11
      P[ 370] <= 9'b110001111; // Load the target box with 15
      P[ 371] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 372] <= 9'b000000000; // Load the constant box with 0
      P[ 373] <= 9'b101001100; // Load the source box with 12
      P[ 374] <= 9'b110001111; // Load the target box with 15
      P[ 375] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 376] <= 9'b000000001; // Load the constant box with 1
      P[ 377] <= 9'b101000000; // Load the source box with 0
      P[ 378] <= 9'b110000000; // Load the target box with 0
      P[ 379] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 380] <= 9'b000000000; // Load the constant box with 0
      P[ 381] <= 9'b101001111; // Load the source box with 15
      P[ 382] <= 9'b110000000; // Load the target box with 0
      P[ 383] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 384] <= 9'b011111010; // Load the constant box with 250
      P[ 385] <= 9'b101000000; // Load the source box with 0
      P[ 386] <= 9'b110000000; // Load the target box with 0
      P[ 387] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 388] <= 9'b000000000; // Load the constant box with 0
      P[ 389] <= 9'b101000000; // Load the source box with 0
      P[ 390] <= 9'b110000001; // Load the target box with 1
      P[ 391] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 392] <= 9'b000000001; // Load the constant box with 1
      P[ 393] <= 9'b101000000; // Load the source box with 0
      P[ 394] <= 9'b110000000; // Load the target box with 0
      P[ 395] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 396] <= 9'b000000000; // Load the constant box with 0
      P[ 397] <= 9'b101000000; // Load the source box with 0
      P[ 398] <= 9'b110001110; // Load the target box with 14
      P[ 399] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 400] <= 9'b000000000; // Load the constant box with 0
      P[ 401] <= 9'b101000010; // Load the source box with 2
      P[ 402] <= 9'b110000001; // Load the target box with 1
      P[ 403] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 404] <= 9'b000000000; // Load the constant box with 0
      P[ 405] <= 9'b101000011; // Load the source box with 3
      P[ 406] <= 9'b110000001; // Load the target box with 1
      P[ 407] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 408] <= 9'b000000000; // Load the constant box with 0
      P[ 409] <= 9'b101000100; // Load the source box with 4
      P[ 410] <= 9'b110000001; // Load the target box with 1
      P[ 411] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 412] <= 9'b000000000; // Load the constant box with 0
      P[ 413] <= 9'b101000101; // Load the source box with 5
      P[ 414] <= 9'b110000001; // Load the target box with 1
      P[ 415] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 416] <= 9'b000000000; // Load the constant box with 0
      P[ 417] <= 9'b101000110; // Load the source box with 6
      P[ 418] <= 9'b110000001; // Load the target box with 1
      P[ 419] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 420] <= 9'b000000000; // Load the constant box with 0
      P[ 421] <= 9'b101000111; // Load the source box with 7
      P[ 422] <= 9'b110000001; // Load the target box with 1
      P[ 423] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 424] <= 9'b000000000; // Load the constant box with 0
      P[ 425] <= 9'b101001000; // Load the source box with 8
      P[ 426] <= 9'b110000001; // Load the target box with 1
      P[ 427] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 428] <= 9'b000000000; // Load the constant box with 0
      P[ 429] <= 9'b101001001; // Load the source box with 9
      P[ 430] <= 9'b110000001; // Load the target box with 1
      P[ 431] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 432] <= 9'b000000000; // Load the constant box with 0
      P[ 433] <= 9'b101001010; // Load the source box with 10
      P[ 434] <= 9'b110000001; // Load the target box with 1
      P[ 435] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 436] <= 9'b000000000; // Load the constant box with 0
      P[ 437] <= 9'b101001011; // Load the source box with 11
      P[ 438] <= 9'b110000001; // Load the target box with 1
      P[ 439] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 440] <= 9'b000000000; // Load the constant box with 0
      P[ 441] <= 9'b101001100; // Load the source box with 12
      P[ 442] <= 9'b110000001; // Load the target box with 1
      P[ 443] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 444] <= 9'b000000001; // Load the constant box with 1
      P[ 445] <= 9'b101000000; // Load the source box with 0
      P[ 446] <= 9'b110000000; // Load the target box with 0
      P[ 447] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 448] <= 9'b000000000; // Load the constant box with 0
      P[ 449] <= 9'b101000001; // Load the source box with 1
      P[ 450] <= 9'b110000000; // Load the target box with 0
      P[ 451] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 452] <= 9'b011110110; // Load the constant box with 246
      P[ 453] <= 9'b101000000; // Load the source box with 0
      P[ 454] <= 9'b110000000; // Load the target box with 0
      P[ 455] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 456] <= 9'b000000000; // Load the constant box with 0
      P[ 457] <= 9'b101000000; // Load the source box with 0
      P[ 458] <= 9'b110001110; // Load the target box with 14
      P[ 459] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 460] <= 9'b011111100; // Load the constant box with 252
      P[ 461] <= 9'b101001101; // Load the source box with 13
      P[ 462] <= 9'b110000000; // Load the target box with 0
      P[ 463] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 464] <= 9'b011111011; // Load the constant box with 251
      P[ 465] <= 9'b101001110; // Load the source box with 14
      P[ 466] <= 9'b110000000; // Load the target box with 0
      P[ 467] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 468] <= 9'b000000000; // Load the constant box with 0
      P[ 469] <= 9'b101000000; // Load the source box with 0
      P[ 470] <= 9'b110000000; // Load the target box with 0
      P[ 471] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task automatic load_Program1;                                                 // Program 1 low
    begin
      $display("Program 1");
      P[   0] <= 9'b000011110; // Load the constant box with 30
      P[   1] <= 9'b101000000; // Load the source box with 0
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   4] <= 9'b000000001; // Load the constant box with 1
      P[   5] <= 9'b101000000; // Load the source box with 0
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001001; // label: Create and set a label
      P[   8] <= 9'b000000000; // Load the constant box with 0
      P[   9] <= 9'b101000000; // Load the source box with 0
      P[  10] <= 9'b110000000; // Load the target box with 0
      P[  11] <= 9'b111000101; // dec: Decrement a register by one
      P[  12] <= 9'b000000000; // Load the constant box with 0
      P[  13] <= 9'b101000000; // Load the source box with 0
      P[  14] <= 9'b110000001; // Load the target box with 1
      P[  15] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[  16] <= 9'b000000000; // Load the constant box with 0
      P[  17] <= 9'b101000000; // Load the source box with 0
      P[  18] <= 9'b110000000; // Load the target box with 0
      P[  19] <= 9'b111000101; // dec: Decrement a register by one
      P[  20] <= 9'b000000000; // Load the constant box with 0
      P[  21] <= 9'b101000000; // Load the source box with 0
      P[  22] <= 9'b110000010; // Load the target box with 2
      P[  23] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[  24] <= 9'b011111111; // Load the constant box with 255
      P[  25] <= 9'b101000000; // Load the source box with 0
      P[  26] <= 9'b110000000; // Load the target box with 0
      P[  27] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  28] <= 9'b011111110; // Load the constant box with 254
      P[  29] <= 9'b101000001; // Load the source box with 1
      P[  30] <= 9'b110000000; // Load the target box with 0
      P[  31] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  32] <= 9'b011111101; // Load the constant box with 253
      P[  33] <= 9'b101000010; // Load the source box with 2
      P[  34] <= 9'b110000000; // Load the target box with 0
      P[  35] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  36] <= 9'b011111110; // Load the constant box with 254
      P[  37] <= 9'b101000001; // Load the source box with 1
      P[  38] <= 9'b110000000; // Load the target box with 0
      P[  39] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[  40] <= 9'b011111101; // Load the constant box with 253
      P[  41] <= 9'b101000010; // Load the source box with 2
      P[  42] <= 9'b110000000; // Load the target box with 0
      P[  43] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[  44] <= 9'b000001000; // Load the constant box with 8
      P[  45] <= 9'b101000001; // Load the source box with 1
      P[  46] <= 9'b110000000; // Load the target box with 0
      P[  47] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  48] <= 9'b000000000; // Load the constant box with 0
      P[  49] <= 9'b101000010; // Load the source box with 2
      P[  50] <= 9'b110000001; // Load the target box with 1
      P[  51] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[  52] <= 9'b000000000; // Load the constant box with 0
      P[  53] <= 9'b101000001; // Load the source box with 1
      P[  54] <= 9'b110000010; // Load the target box with 2
      P[  55] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  56] <= 9'b000000101; // Load the constant box with 5
      P[  57] <= 9'b101000010; // Load the source box with 2
      P[  58] <= 9'b110000000; // Load the target box with 0
      P[  59] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  60] <= 9'b000001111; // Load the constant box with 15
      P[  61] <= 9'b101000010; // Load the source box with 2
      P[  62] <= 9'b110000000; // Load the target box with 0
      P[  63] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  64] <= 9'b000000000; // Load the constant box with 0
      P[  65] <= 9'b101000001; // Load the source box with 1
      P[  66] <= 9'b110000011; // Load the target box with 3
      P[  67] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  68] <= 9'b000000110; // Load the constant box with 6
      P[  69] <= 9'b101000011; // Load the source box with 3
      P[  70] <= 9'b110000000; // Load the target box with 0
      P[  71] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  72] <= 9'b000001111; // Load the constant box with 15
      P[  73] <= 9'b101000011; // Load the source box with 3
      P[  74] <= 9'b110000000; // Load the target box with 0
      P[  75] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  76] <= 9'b000000000; // Load the constant box with 0
      P[  77] <= 9'b101000001; // Load the source box with 1
      P[  78] <= 9'b110000100; // Load the target box with 4
      P[  79] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  80] <= 9'b000000111; // Load the constant box with 7
      P[  81] <= 9'b101000100; // Load the source box with 4
      P[  82] <= 9'b110000000; // Load the target box with 0
      P[  83] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  84] <= 9'b000001111; // Load the constant box with 15
      P[  85] <= 9'b101000100; // Load the source box with 4
      P[  86] <= 9'b110000000; // Load the target box with 0
      P[  87] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  88] <= 9'b000000000; // Load the constant box with 0
      P[  89] <= 9'b101000001; // Load the source box with 1
      P[  90] <= 9'b110000101; // Load the target box with 5
      P[  91] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  92] <= 9'b000001000; // Load the constant box with 8
      P[  93] <= 9'b101000101; // Load the source box with 5
      P[  94] <= 9'b110000000; // Load the target box with 0
      P[  95] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  96] <= 9'b000001111; // Load the constant box with 15
      P[  97] <= 9'b101000101; // Load the source box with 5
      P[  98] <= 9'b110000000; // Load the target box with 0
      P[  99] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 100] <= 9'b000000000; // Load the constant box with 0
      P[ 101] <= 9'b101000001; // Load the source box with 1
      P[ 102] <= 9'b110000110; // Load the target box with 6
      P[ 103] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 104] <= 9'b000001001; // Load the constant box with 9
      P[ 105] <= 9'b101000110; // Load the source box with 6
      P[ 106] <= 9'b110000000; // Load the target box with 0
      P[ 107] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 108] <= 9'b000001111; // Load the constant box with 15
      P[ 109] <= 9'b101000110; // Load the source box with 6
      P[ 110] <= 9'b110000000; // Load the target box with 0
      P[ 111] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 112] <= 9'b000000000; // Load the constant box with 0
      P[ 113] <= 9'b101000001; // Load the source box with 1
      P[ 114] <= 9'b110000111; // Load the target box with 7
      P[ 115] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 116] <= 9'b000001010; // Load the constant box with 10
      P[ 117] <= 9'b101000111; // Load the source box with 7
      P[ 118] <= 9'b110000000; // Load the target box with 0
      P[ 119] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 120] <= 9'b000001111; // Load the constant box with 15
      P[ 121] <= 9'b101000111; // Load the source box with 7
      P[ 122] <= 9'b110000000; // Load the target box with 0
      P[ 123] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 124] <= 9'b000000000; // Load the constant box with 0
      P[ 125] <= 9'b101000001; // Load the source box with 1
      P[ 126] <= 9'b110001000; // Load the target box with 8
      P[ 127] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 128] <= 9'b000001011; // Load the constant box with 11
      P[ 129] <= 9'b101001000; // Load the source box with 8
      P[ 130] <= 9'b110000000; // Load the target box with 0
      P[ 131] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 132] <= 9'b000001111; // Load the constant box with 15
      P[ 133] <= 9'b101001000; // Load the source box with 8
      P[ 134] <= 9'b110000000; // Load the target box with 0
      P[ 135] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 136] <= 9'b000000000; // Load the constant box with 0
      P[ 137] <= 9'b101000001; // Load the source box with 1
      P[ 138] <= 9'b110001001; // Load the target box with 9
      P[ 139] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 140] <= 9'b000001100; // Load the constant box with 12
      P[ 141] <= 9'b101001001; // Load the source box with 9
      P[ 142] <= 9'b110000000; // Load the target box with 0
      P[ 143] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 144] <= 9'b000001111; // Load the constant box with 15
      P[ 145] <= 9'b101001001; // Load the source box with 9
      P[ 146] <= 9'b110000000; // Load the target box with 0
      P[ 147] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 148] <= 9'b000000000; // Load the constant box with 0
      P[ 149] <= 9'b101000001; // Load the source box with 1
      P[ 150] <= 9'b110001010; // Load the target box with 10
      P[ 151] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 152] <= 9'b000001101; // Load the constant box with 13
      P[ 153] <= 9'b101001010; // Load the source box with 10
      P[ 154] <= 9'b110000000; // Load the target box with 0
      P[ 155] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 156] <= 9'b000001111; // Load the constant box with 15
      P[ 157] <= 9'b101001010; // Load the source box with 10
      P[ 158] <= 9'b110000000; // Load the target box with 0
      P[ 159] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 160] <= 9'b000000000; // Load the constant box with 0
      P[ 161] <= 9'b101000001; // Load the source box with 1
      P[ 162] <= 9'b110001011; // Load the target box with 11
      P[ 163] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 164] <= 9'b000001110; // Load the constant box with 14
      P[ 165] <= 9'b101001011; // Load the source box with 11
      P[ 166] <= 9'b110000000; // Load the target box with 0
      P[ 167] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 168] <= 9'b000001111; // Load the constant box with 15
      P[ 169] <= 9'b101001011; // Load the source box with 11
      P[ 170] <= 9'b110000000; // Load the target box with 0
      P[ 171] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 172] <= 9'b000000000; // Load the constant box with 0
      P[ 173] <= 9'b101000001; // Load the source box with 1
      P[ 174] <= 9'b110001100; // Load the target box with 12
      P[ 175] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 176] <= 9'b000001111; // Load the constant box with 15
      P[ 177] <= 9'b101001100; // Load the source box with 12
      P[ 178] <= 9'b110000000; // Load the target box with 0
      P[ 179] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 180] <= 9'b000001111; // Load the constant box with 15
      P[ 181] <= 9'b101001100; // Load the source box with 12
      P[ 182] <= 9'b110000000; // Load the target box with 0
      P[ 183] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 184] <= 9'b000000000; // Load the constant box with 0
      P[ 185] <= 9'b101000001; // Load the source box with 1
      P[ 186] <= 9'b110001101; // Load the target box with 13
      P[ 187] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 188] <= 9'b000000101; // Load the constant box with 5
      P[ 189] <= 9'b101001101; // Load the source box with 13
      P[ 190] <= 9'b110000000; // Load the target box with 0
      P[ 191] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 192] <= 9'b000001001; // Load the constant box with 9
      P[ 193] <= 9'b101001101; // Load the source box with 13
      P[ 194] <= 9'b110000000; // Load the target box with 0
      P[ 195] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 196] <= 9'b000000001; // Load the constant box with 1
      P[ 197] <= 9'b101001101; // Load the source box with 13
      P[ 198] <= 9'b110000000; // Load the target box with 0
      P[ 199] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 200] <= 9'b000000000; // Load the constant box with 0
      P[ 201] <= 9'b101000001; // Load the source box with 1
      P[ 202] <= 9'b110001110; // Load the target box with 14
      P[ 203] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 204] <= 9'b000001000; // Load the constant box with 8
      P[ 205] <= 9'b101001110; // Load the source box with 14
      P[ 206] <= 9'b110000000; // Load the target box with 0
      P[ 207] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 208] <= 9'b000001101; // Load the constant box with 13
      P[ 209] <= 9'b101001110; // Load the source box with 14
      P[ 210] <= 9'b110000000; // Load the target box with 0
      P[ 211] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 212] <= 9'b000000101; // Load the constant box with 5
      P[ 213] <= 9'b101001110; // Load the source box with 14
      P[ 214] <= 9'b110000000; // Load the target box with 0
      P[ 215] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 216] <= 9'b000000000; // Load the constant box with 0
      P[ 217] <= 9'b101000001; // Load the source box with 1
      P[ 218] <= 9'b110001111; // Load the target box with 15
      P[ 219] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 220] <= 9'b000001111; // Load the constant box with 15
      P[ 221] <= 9'b101001111; // Load the source box with 15
      P[ 222] <= 9'b110000000; // Load the target box with 0
      P[ 223] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 224] <= 9'b000001100; // Load the constant box with 12
      P[ 225] <= 9'b101001111; // Load the source box with 15
      P[ 226] <= 9'b110000000; // Load the target box with 0
      P[ 227] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 228] <= 9'b000000000; // Load the constant box with 0
      P[ 229] <= 9'b101001111; // Load the source box with 15
      P[ 230] <= 9'b110001110; // Load the target box with 14
      P[ 231] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 232] <= 9'b000000000; // Load the constant box with 0
      P[ 233] <= 9'b101000010; // Load the source box with 2
      P[ 234] <= 9'b110001111; // Load the target box with 15
      P[ 235] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 236] <= 9'b000000000; // Load the constant box with 0
      P[ 237] <= 9'b101000011; // Load the source box with 3
      P[ 238] <= 9'b110001111; // Load the target box with 15
      P[ 239] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 240] <= 9'b000000000; // Load the constant box with 0
      P[ 241] <= 9'b101000100; // Load the source box with 4
      P[ 242] <= 9'b110001111; // Load the target box with 15
      P[ 243] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 244] <= 9'b000000000; // Load the constant box with 0
      P[ 245] <= 9'b101000101; // Load the source box with 5
      P[ 246] <= 9'b110001111; // Load the target box with 15
      P[ 247] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 248] <= 9'b000000000; // Load the constant box with 0
      P[ 249] <= 9'b101000110; // Load the source box with 6
      P[ 250] <= 9'b110001111; // Load the target box with 15
      P[ 251] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 252] <= 9'b000000000; // Load the constant box with 0
      P[ 253] <= 9'b101000111; // Load the source box with 7
      P[ 254] <= 9'b110001111; // Load the target box with 15
      P[ 255] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 256] <= 9'b000000000; // Load the constant box with 0
      P[ 257] <= 9'b101001000; // Load the source box with 8
      P[ 258] <= 9'b110001111; // Load the target box with 15
      P[ 259] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 260] <= 9'b000000001; // Load the constant box with 1
      P[ 261] <= 9'b101000000; // Load the source box with 0
      P[ 262] <= 9'b110000000; // Load the target box with 0
      P[ 263] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 264] <= 9'b000000000; // Load the constant box with 0
      P[ 265] <= 9'b101001111; // Load the source box with 15
      P[ 266] <= 9'b110000000; // Load the target box with 0
      P[ 267] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 268] <= 9'b011110111; // Load the constant box with 247
      P[ 269] <= 9'b101000000; // Load the source box with 0
      P[ 270] <= 9'b110000000; // Load the target box with 0
      P[ 271] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 272] <= 9'b000000000; // Load the constant box with 0
      P[ 273] <= 9'b101000000; // Load the source box with 0
      P[ 274] <= 9'b110000001; // Load the target box with 1
      P[ 275] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 276] <= 9'b000000000; // Load the constant box with 0
      P[ 277] <= 9'b101000000; // Load the source box with 0
      P[ 278] <= 9'b110001101; // Load the target box with 13
      P[ 279] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 280] <= 9'b000000000; // Load the constant box with 0
      P[ 281] <= 9'b101000010; // Load the source box with 2
      P[ 282] <= 9'b110001111; // Load the target box with 15
      P[ 283] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 284] <= 9'b000000000; // Load the constant box with 0
      P[ 285] <= 9'b101000011; // Load the source box with 3
      P[ 286] <= 9'b110001111; // Load the target box with 15
      P[ 287] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 288] <= 9'b000000000; // Load the constant box with 0
      P[ 289] <= 9'b101000100; // Load the source box with 4
      P[ 290] <= 9'b110001111; // Load the target box with 15
      P[ 291] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 292] <= 9'b000000000; // Load the constant box with 0
      P[ 293] <= 9'b101000101; // Load the source box with 5
      P[ 294] <= 9'b110001111; // Load the target box with 15
      P[ 295] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 296] <= 9'b000000000; // Load the constant box with 0
      P[ 297] <= 9'b101001001; // Load the source box with 9
      P[ 298] <= 9'b110001111; // Load the target box with 15
      P[ 299] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 300] <= 9'b000000000; // Load the constant box with 0
      P[ 301] <= 9'b101001010; // Load the source box with 10
      P[ 302] <= 9'b110001111; // Load the target box with 15
      P[ 303] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 304] <= 9'b000000000; // Load the constant box with 0
      P[ 305] <= 9'b101001011; // Load the source box with 11
      P[ 306] <= 9'b110001111; // Load the target box with 15
      P[ 307] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 308] <= 9'b000000001; // Load the constant box with 1
      P[ 309] <= 9'b101000000; // Load the source box with 0
      P[ 310] <= 9'b110000000; // Load the target box with 0
      P[ 311] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 312] <= 9'b000000000; // Load the constant box with 0
      P[ 313] <= 9'b101001111; // Load the source box with 15
      P[ 314] <= 9'b110000000; // Load the target box with 0
      P[ 315] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 316] <= 9'b011111000; // Load the constant box with 248
      P[ 317] <= 9'b101000000; // Load the source box with 0
      P[ 318] <= 9'b110000000; // Load the target box with 0
      P[ 319] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 320] <= 9'b000000000; // Load the constant box with 0
      P[ 321] <= 9'b101000000; // Load the source box with 0
      P[ 322] <= 9'b110000001; // Load the target box with 1
      P[ 323] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 324] <= 9'b000000100; // Load the constant box with 4
      P[ 325] <= 9'b101000000; // Load the source box with 0
      P[ 326] <= 9'b110000000; // Load the target box with 0
      P[ 327] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 328] <= 9'b000000000; // Load the constant box with 0
      P[ 329] <= 9'b101000000; // Load the source box with 0
      P[ 330] <= 9'b110001110; // Load the target box with 14
      P[ 331] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 332] <= 9'b000000000; // Load the constant box with 0
      P[ 333] <= 9'b101000010; // Load the source box with 2
      P[ 334] <= 9'b110001111; // Load the target box with 15
      P[ 335] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 336] <= 9'b000000000; // Load the constant box with 0
      P[ 337] <= 9'b101000011; // Load the source box with 3
      P[ 338] <= 9'b110001111; // Load the target box with 15
      P[ 339] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 340] <= 9'b000000000; // Load the constant box with 0
      P[ 341] <= 9'b101000110; // Load the source box with 6
      P[ 342] <= 9'b110001111; // Load the target box with 15
      P[ 343] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 344] <= 9'b000000000; // Load the constant box with 0
      P[ 345] <= 9'b101000111; // Load the source box with 7
      P[ 346] <= 9'b110001111; // Load the target box with 15
      P[ 347] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 348] <= 9'b000000000; // Load the constant box with 0
      P[ 349] <= 9'b101001001; // Load the source box with 9
      P[ 350] <= 9'b110001111; // Load the target box with 15
      P[ 351] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 352] <= 9'b000000000; // Load the constant box with 0
      P[ 353] <= 9'b101001010; // Load the source box with 10
      P[ 354] <= 9'b110001111; // Load the target box with 15
      P[ 355] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 356] <= 9'b000000000; // Load the constant box with 0
      P[ 357] <= 9'b101001100; // Load the source box with 12
      P[ 358] <= 9'b110001111; // Load the target box with 15
      P[ 359] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 360] <= 9'b000000001; // Load the constant box with 1
      P[ 361] <= 9'b101000000; // Load the source box with 0
      P[ 362] <= 9'b110000000; // Load the target box with 0
      P[ 363] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 364] <= 9'b000000000; // Load the constant box with 0
      P[ 365] <= 9'b101001111; // Load the source box with 15
      P[ 366] <= 9'b110000000; // Load the target box with 0
      P[ 367] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 368] <= 9'b011111001; // Load the constant box with 249
      P[ 369] <= 9'b101000000; // Load the source box with 0
      P[ 370] <= 9'b110000000; // Load the target box with 0
      P[ 371] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 372] <= 9'b000000000; // Load the constant box with 0
      P[ 373] <= 9'b101000000; // Load the source box with 0
      P[ 374] <= 9'b110000001; // Load the target box with 1
      P[ 375] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 376] <= 9'b000000010; // Load the constant box with 2
      P[ 377] <= 9'b101000000; // Load the source box with 0
      P[ 378] <= 9'b110000000; // Load the target box with 0
      P[ 379] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 380] <= 9'b000000000; // Load the constant box with 0
      P[ 381] <= 9'b101000000; // Load the source box with 0
      P[ 382] <= 9'b110001110; // Load the target box with 14
      P[ 383] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 384] <= 9'b000000000; // Load the constant box with 0
      P[ 385] <= 9'b101000010; // Load the source box with 2
      P[ 386] <= 9'b110001111; // Load the target box with 15
      P[ 387] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 388] <= 9'b000000000; // Load the constant box with 0
      P[ 389] <= 9'b101000100; // Load the source box with 4
      P[ 390] <= 9'b110001111; // Load the target box with 15
      P[ 391] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 392] <= 9'b000000000; // Load the constant box with 0
      P[ 393] <= 9'b101000110; // Load the source box with 6
      P[ 394] <= 9'b110001111; // Load the target box with 15
      P[ 395] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 396] <= 9'b000000000; // Load the constant box with 0
      P[ 397] <= 9'b101001000; // Load the source box with 8
      P[ 398] <= 9'b110001111; // Load the target box with 15
      P[ 399] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 400] <= 9'b000000000; // Load the constant box with 0
      P[ 401] <= 9'b101001001; // Load the source box with 9
      P[ 402] <= 9'b110001111; // Load the target box with 15
      P[ 403] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 404] <= 9'b000000000; // Load the constant box with 0
      P[ 405] <= 9'b101001011; // Load the source box with 11
      P[ 406] <= 9'b110001111; // Load the target box with 15
      P[ 407] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 408] <= 9'b000000000; // Load the constant box with 0
      P[ 409] <= 9'b101001100; // Load the source box with 12
      P[ 410] <= 9'b110001111; // Load the target box with 15
      P[ 411] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 412] <= 9'b000000001; // Load the constant box with 1
      P[ 413] <= 9'b101000000; // Load the source box with 0
      P[ 414] <= 9'b110000000; // Load the target box with 0
      P[ 415] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 416] <= 9'b000000000; // Load the constant box with 0
      P[ 417] <= 9'b101001111; // Load the source box with 15
      P[ 418] <= 9'b110000000; // Load the target box with 0
      P[ 419] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 420] <= 9'b011111010; // Load the constant box with 250
      P[ 421] <= 9'b101000000; // Load the source box with 0
      P[ 422] <= 9'b110000000; // Load the target box with 0
      P[ 423] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 424] <= 9'b000000000; // Load the constant box with 0
      P[ 425] <= 9'b101000000; // Load the source box with 0
      P[ 426] <= 9'b110000001; // Load the target box with 1
      P[ 427] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 428] <= 9'b000000001; // Load the constant box with 1
      P[ 429] <= 9'b101000000; // Load the source box with 0
      P[ 430] <= 9'b110000000; // Load the target box with 0
      P[ 431] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 432] <= 9'b000000000; // Load the constant box with 0
      P[ 433] <= 9'b101000000; // Load the source box with 0
      P[ 434] <= 9'b110001110; // Load the target box with 14
      P[ 435] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 436] <= 9'b000000000; // Load the constant box with 0
      P[ 437] <= 9'b101000010; // Load the source box with 2
      P[ 438] <= 9'b110000001; // Load the target box with 1
      P[ 439] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 440] <= 9'b000000000; // Load the constant box with 0
      P[ 441] <= 9'b101000011; // Load the source box with 3
      P[ 442] <= 9'b110000001; // Load the target box with 1
      P[ 443] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 444] <= 9'b000000000; // Load the constant box with 0
      P[ 445] <= 9'b101000100; // Load the source box with 4
      P[ 446] <= 9'b110000001; // Load the target box with 1
      P[ 447] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 448] <= 9'b000000000; // Load the constant box with 0
      P[ 449] <= 9'b101000101; // Load the source box with 5
      P[ 450] <= 9'b110000001; // Load the target box with 1
      P[ 451] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 452] <= 9'b000000000; // Load the constant box with 0
      P[ 453] <= 9'b101000110; // Load the source box with 6
      P[ 454] <= 9'b110000001; // Load the target box with 1
      P[ 455] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 456] <= 9'b000000000; // Load the constant box with 0
      P[ 457] <= 9'b101000111; // Load the source box with 7
      P[ 458] <= 9'b110000001; // Load the target box with 1
      P[ 459] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 460] <= 9'b000000000; // Load the constant box with 0
      P[ 461] <= 9'b101001000; // Load the source box with 8
      P[ 462] <= 9'b110000001; // Load the target box with 1
      P[ 463] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 464] <= 9'b000000000; // Load the constant box with 0
      P[ 465] <= 9'b101001001; // Load the source box with 9
      P[ 466] <= 9'b110000001; // Load the target box with 1
      P[ 467] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 468] <= 9'b000000000; // Load the constant box with 0
      P[ 469] <= 9'b101001010; // Load the source box with 10
      P[ 470] <= 9'b110000001; // Load the target box with 1
      P[ 471] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 472] <= 9'b000000000; // Load the constant box with 0
      P[ 473] <= 9'b101001011; // Load the source box with 11
      P[ 474] <= 9'b110000001; // Load the target box with 1
      P[ 475] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 476] <= 9'b000000000; // Load the constant box with 0
      P[ 477] <= 9'b101001100; // Load the source box with 12
      P[ 478] <= 9'b110000001; // Load the target box with 1
      P[ 479] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 480] <= 9'b000000001; // Load the constant box with 1
      P[ 481] <= 9'b101000000; // Load the source box with 0
      P[ 482] <= 9'b110000000; // Load the target box with 0
      P[ 483] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 484] <= 9'b000000000; // Load the constant box with 0
      P[ 485] <= 9'b101000001; // Load the source box with 1
      P[ 486] <= 9'b110000000; // Load the target box with 0
      P[ 487] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 488] <= 9'b011110110; // Load the constant box with 246
      P[ 489] <= 9'b101000000; // Load the source box with 0
      P[ 490] <= 9'b110000000; // Load the target box with 0
      P[ 491] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 492] <= 9'b000000000; // Load the constant box with 0
      P[ 493] <= 9'b101000000; // Load the source box with 0
      P[ 494] <= 9'b110001110; // Load the target box with 14
      P[ 495] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 496] <= 9'b011111100; // Load the constant box with 252
      P[ 497] <= 9'b101001101; // Load the source box with 13
      P[ 498] <= 9'b110000000; // Load the target box with 0
      P[ 499] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 500] <= 9'b011111011; // Load the constant box with 251
      P[ 501] <= 9'b101001110; // Load the source box with 14
      P[ 502] <= 9'b110000000; // Load the target box with 0
      P[ 503] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 504] <= 9'b011111111; // Load the constant box with 255
      P[ 505] <= 9'b101000000; // Load the source box with 0
      P[ 506] <= 9'b110000000; // Load the target box with 0
      P[ 507] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 508] <= 9'b011111100; // Load the constant box with 252
      P[ 509] <= 9'b101001101; // Load the source box with 13
      P[ 510] <= 9'b110000000; // Load the target box with 0
      P[ 511] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 512] <= 9'b011111011; // Load the constant box with 251
      P[ 513] <= 9'b101001110; // Load the source box with 14
      P[ 514] <= 9'b110000000; // Load the target box with 0
      P[ 515] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 516] <= 9'b000011110; // Load the constant box with 30
      P[ 517] <= 9'b101000001; // Load the source box with 1
      P[ 518] <= 9'b110000000; // Load the target box with 0
      P[ 519] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 520] <= 9'b000000000; // Load the constant box with 0
      P[ 521] <= 9'b101000000; // Load the source box with 0
      P[ 522] <= 9'b110000001; // Load the target box with 1
      P[ 523] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 524] <= 9'b000000000; // Load the constant box with 0
      P[ 525] <= 9'b101000001; // Load the source box with 1
      P[ 526] <= 9'b110001110; // Load the target box with 14
      P[ 527] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[ 528] <= 9'b000000000; // Load the constant box with 0
      P[ 529] <= 9'b101000001; // Load the source box with 1
      P[ 530] <= 9'b110000000; // Load the target box with 0
      P[ 531] <= 9'b111000110; // inc: Increment a register by one
      P[ 532] <= 9'b000000000; // Load the constant box with 0
      P[ 533] <= 9'b101000001; // Load the source box with 1
      P[ 534] <= 9'b110001101; // Load the target box with 13
      P[ 535] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[ 536] <= 9'b000000001; // Load the constant box with 1
      P[ 537] <= 9'b101000000; // Load the source box with 0
      P[ 538] <= 9'b110000000; // Load the target box with 0
      P[ 539] <= 9'b111000111; // jumpIfNotZero: Jump backwards to the specified location in the program if the register is not zero - useful for constructing for loops
      P[ 540] <= 9'b000000000; // Load the constant box with 0
      P[ 541] <= 9'b101000000; // Load the source box with 0
      P[ 542] <= 9'b110000000; // Load the target box with 0
      P[ 543] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task automatic load_Program2;                                                           // Program 2
    begin
      $display("Program 2");
      P[   0] <= 9'b001011110; // Load the constant box with 94
      P[   1] <= 9'b101000000; // Load the source box with 0
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   4] <= 9'b000001101; // Load the constant box with 13
      P[   5] <= 9'b101000000; // Load the source box with 0
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001001; // label: Create and set a label
      P[   8] <= 9'b000000000; // Load the constant box with 0
      P[   9] <= 9'b101000000; // Load the source box with 0
      P[  10] <= 9'b110000000; // Load the target box with 0
      P[  11] <= 9'b111000101; // dec: Decrement a register by one
      P[  12] <= 9'b000000000; // Load the constant box with 0
      P[  13] <= 9'b101000000; // Load the source box with 0
      P[  14] <= 9'b110000010; // Load the target box with 2
      P[  15] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[  16] <= 9'b000000000; // Load the constant box with 0
      P[  17] <= 9'b101000000; // Load the source box with 0
      P[  18] <= 9'b110000000; // Load the target box with 0
      P[  19] <= 9'b111000101; // dec: Decrement a register by one
      P[  20] <= 9'b000000000; // Load the constant box with 0
      P[  21] <= 9'b101000000; // Load the source box with 0
      P[  22] <= 9'b110000001; // Load the target box with 1
      P[  23] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[  24] <= 9'b000000000; // Load the constant box with 0
      P[  25] <= 9'b101000010; // Load the source box with 2
      P[  26] <= 9'b110000011; // Load the target box with 3
      P[  27] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  28] <= 9'b000000101; // Load the constant box with 5
      P[  29] <= 9'b101000011; // Load the source box with 3
      P[  30] <= 9'b110000000; // Load the target box with 0
      P[  31] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  32] <= 9'b000000000; // Load the constant box with 0
      P[  33] <= 9'b101000010; // Load the source box with 2
      P[  34] <= 9'b110000100; // Load the target box with 4
      P[  35] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  36] <= 9'b000000001; // Load the constant box with 1
      P[  37] <= 9'b101000100; // Load the source box with 4
      P[  38] <= 9'b110000000; // Load the target box with 0
      P[  39] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  40] <= 9'b000001100; // Load the constant box with 12
      P[  41] <= 9'b101000100; // Load the source box with 4
      P[  42] <= 9'b110000000; // Load the target box with 0
      P[  43] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  44] <= 9'b000001000; // Load the constant box with 8
      P[  45] <= 9'b101000100; // Load the source box with 4
      P[  46] <= 9'b110000000; // Load the target box with 0
      P[  47] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  48] <= 9'b000000000; // Load the constant box with 0
      P[  49] <= 9'b101000001; // Load the source box with 1
      P[  50] <= 9'b110000101; // Load the target box with 5
      P[  51] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  52] <= 9'b000000101; // Load the constant box with 5
      P[  53] <= 9'b101000101; // Load the source box with 5
      P[  54] <= 9'b110000000; // Load the target box with 0
      P[  55] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  56] <= 9'b000000001; // Load the constant box with 1
      P[  57] <= 9'b101000101; // Load the source box with 5
      P[  58] <= 9'b110000000; // Load the target box with 0
      P[  59] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  60] <= 9'b000000000; // Load the constant box with 0
      P[  61] <= 9'b101000101; // Load the source box with 5
      P[  62] <= 9'b110000100; // Load the target box with 4
      P[  63] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[  64] <= 9'b000000000; // Load the constant box with 0
      P[  65] <= 9'b101000001; // Load the source box with 1
      P[  66] <= 9'b110000101; // Load the target box with 5
      P[  67] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  68] <= 9'b000001100; // Load the constant box with 12
      P[  69] <= 9'b101000101; // Load the source box with 5
      P[  70] <= 9'b110000000; // Load the target box with 0
      P[  71] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  72] <= 9'b000001111; // Load the constant box with 15
      P[  73] <= 9'b101000101; // Load the source box with 5
      P[  74] <= 9'b110000000; // Load the target box with 0
      P[  75] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  76] <= 9'b000000000; // Load the constant box with 0
      P[  77] <= 9'b101000101; // Load the source box with 5
      P[  78] <= 9'b110000100; // Load the target box with 4
      P[  79] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[  80] <= 9'b011111111; // Load the constant box with 255
      P[  81] <= 9'b101000000; // Load the source box with 0
      P[  82] <= 9'b110000000; // Load the target box with 0
      P[  83] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  84] <= 9'b011111110; // Load the constant box with 254
      P[  85] <= 9'b101000011; // Load the source box with 3
      P[  86] <= 9'b110000000; // Load the target box with 0
      P[  87] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  88] <= 9'b011111101; // Load the constant box with 253
      P[  89] <= 9'b101000100; // Load the source box with 4
      P[  90] <= 9'b110000000; // Load the target box with 0
      P[  91] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[  92] <= 9'b000000000; // Load the constant box with 0
      P[  93] <= 9'b101000010; // Load the source box with 2
      P[  94] <= 9'b110000011; // Load the target box with 3
      P[  95] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  96] <= 9'b000000001; // Load the constant box with 1
      P[  97] <= 9'b101000100; // Load the source box with 4
      P[  98] <= 9'b110000000; // Load the target box with 0
      P[  99] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 100] <= 9'b000000000; // Load the constant box with 0
      P[ 101] <= 9'b101000011; // Load the source box with 3
      P[ 102] <= 9'b110000100; // Load the target box with 4
      P[ 103] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 104] <= 9'b011110010; // Load the constant box with 242
      P[ 105] <= 9'b101000100; // Load the source box with 4
      P[ 106] <= 9'b110000000; // Load the target box with 0
      P[ 107] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 108] <= 9'b000000000; // Load the constant box with 0
      P[ 109] <= 9'b101000001; // Load the source box with 1
      P[ 110] <= 9'b110000011; // Load the target box with 3
      P[ 111] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 112] <= 9'b000000100; // Load the constant box with 4
      P[ 113] <= 9'b101000011; // Load the source box with 3
      P[ 114] <= 9'b110000000; // Load the target box with 0
      P[ 115] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 116] <= 9'b000000001; // Load the constant box with 1
      P[ 117] <= 9'b101000100; // Load the source box with 4
      P[ 118] <= 9'b110000000; // Load the target box with 0
      P[ 119] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 120] <= 9'b000000000; // Load the constant box with 0
      P[ 121] <= 9'b101000011; // Load the source box with 3
      P[ 122] <= 9'b110000100; // Load the target box with 4
      P[ 123] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 124] <= 9'b011110011; // Load the constant box with 243
      P[ 125] <= 9'b101000100; // Load the source box with 4
      P[ 126] <= 9'b110000000; // Load the target box with 0
      P[ 127] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 128] <= 9'b000000000; // Load the constant box with 0
      P[ 129] <= 9'b101000001; // Load the source box with 1
      P[ 130] <= 9'b110000011; // Load the target box with 3
      P[ 131] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 132] <= 9'b000000010; // Load the constant box with 2
      P[ 133] <= 9'b101000011; // Load the source box with 3
      P[ 134] <= 9'b110000000; // Load the target box with 0
      P[ 135] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 136] <= 9'b000000001; // Load the constant box with 1
      P[ 137] <= 9'b101000100; // Load the source box with 4
      P[ 138] <= 9'b110000000; // Load the target box with 0
      P[ 139] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 140] <= 9'b000000000; // Load the constant box with 0
      P[ 141] <= 9'b101000011; // Load the source box with 3
      P[ 142] <= 9'b110000100; // Load the target box with 4
      P[ 143] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 144] <= 9'b011110100; // Load the constant box with 244
      P[ 145] <= 9'b101000100; // Load the source box with 4
      P[ 146] <= 9'b110000000; // Load the target box with 0
      P[ 147] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 148] <= 9'b000000000; // Load the constant box with 0
      P[ 149] <= 9'b101000001; // Load the source box with 1
      P[ 150] <= 9'b110000011; // Load the target box with 3
      P[ 151] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 152] <= 9'b000000001; // Load the constant box with 1
      P[ 153] <= 9'b101000011; // Load the source box with 3
      P[ 154] <= 9'b110000000; // Load the target box with 0
      P[ 155] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 156] <= 9'b000000001; // Load the constant box with 1
      P[ 157] <= 9'b101000100; // Load the source box with 4
      P[ 158] <= 9'b110000000; // Load the target box with 0
      P[ 159] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 160] <= 9'b000000000; // Load the constant box with 0
      P[ 161] <= 9'b101000011; // Load the source box with 3
      P[ 162] <= 9'b110000100; // Load the target box with 4
      P[ 163] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 164] <= 9'b011110101; // Load the constant box with 245
      P[ 165] <= 9'b101000100; // Load the source box with 4
      P[ 166] <= 9'b110000000; // Load the target box with 0
      P[ 167] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 168] <= 9'b000000000; // Load the constant box with 0
      P[ 169] <= 9'b101000001; // Load the source box with 1
      P[ 170] <= 9'b110000011; // Load the target box with 3
      P[ 171] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 172] <= 9'b000000001; // Load the constant box with 1
      P[ 173] <= 9'b101000100; // Load the source box with 4
      P[ 174] <= 9'b110000000; // Load the target box with 0
      P[ 175] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 176] <= 9'b000000000; // Load the constant box with 0
      P[ 177] <= 9'b101000011; // Load the source box with 3
      P[ 178] <= 9'b110000100; // Load the target box with 4
      P[ 179] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 180] <= 9'b011110001; // Load the constant box with 241
      P[ 181] <= 9'b101000100; // Load the source box with 4
      P[ 182] <= 9'b110000000; // Load the target box with 0
      P[ 183] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 184] <= 9'b011111110; // Load the constant box with 254
      P[ 185] <= 9'b101000001; // Load the source box with 1
      P[ 186] <= 9'b110000000; // Load the target box with 0
      P[ 187] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 188] <= 9'b011111101; // Load the constant box with 253
      P[ 189] <= 9'b101000010; // Load the source box with 2
      P[ 190] <= 9'b110000000; // Load the target box with 0
      P[ 191] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 192] <= 9'b000001000; // Load the constant box with 8
      P[ 193] <= 9'b101000001; // Load the source box with 1
      P[ 194] <= 9'b110000000; // Load the target box with 0
      P[ 195] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 196] <= 9'b000000000; // Load the constant box with 0
      P[ 197] <= 9'b101000010; // Load the source box with 2
      P[ 198] <= 9'b110000001; // Load the target box with 1
      P[ 199] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 200] <= 9'b000000000; // Load the constant box with 0
      P[ 201] <= 9'b101000001; // Load the source box with 1
      P[ 202] <= 9'b110000010; // Load the target box with 2
      P[ 203] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 204] <= 9'b000000101; // Load the constant box with 5
      P[ 205] <= 9'b101000010; // Load the source box with 2
      P[ 206] <= 9'b110000000; // Load the target box with 0
      P[ 207] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 208] <= 9'b000001111; // Load the constant box with 15
      P[ 209] <= 9'b101000010; // Load the source box with 2
      P[ 210] <= 9'b110000000; // Load the target box with 0
      P[ 211] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 212] <= 9'b000000000; // Load the constant box with 0
      P[ 213] <= 9'b101000001; // Load the source box with 1
      P[ 214] <= 9'b110000011; // Load the target box with 3
      P[ 215] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 216] <= 9'b000000110; // Load the constant box with 6
      P[ 217] <= 9'b101000011; // Load the source box with 3
      P[ 218] <= 9'b110000000; // Load the target box with 0
      P[ 219] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 220] <= 9'b000001111; // Load the constant box with 15
      P[ 221] <= 9'b101000011; // Load the source box with 3
      P[ 222] <= 9'b110000000; // Load the target box with 0
      P[ 223] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 224] <= 9'b000000000; // Load the constant box with 0
      P[ 225] <= 9'b101000001; // Load the source box with 1
      P[ 226] <= 9'b110000100; // Load the target box with 4
      P[ 227] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 228] <= 9'b000000111; // Load the constant box with 7
      P[ 229] <= 9'b101000100; // Load the source box with 4
      P[ 230] <= 9'b110000000; // Load the target box with 0
      P[ 231] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 232] <= 9'b000001111; // Load the constant box with 15
      P[ 233] <= 9'b101000100; // Load the source box with 4
      P[ 234] <= 9'b110000000; // Load the target box with 0
      P[ 235] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 236] <= 9'b000000000; // Load the constant box with 0
      P[ 237] <= 9'b101000001; // Load the source box with 1
      P[ 238] <= 9'b110000101; // Load the target box with 5
      P[ 239] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 240] <= 9'b000001000; // Load the constant box with 8
      P[ 241] <= 9'b101000101; // Load the source box with 5
      P[ 242] <= 9'b110000000; // Load the target box with 0
      P[ 243] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 244] <= 9'b000001111; // Load the constant box with 15
      P[ 245] <= 9'b101000101; // Load the source box with 5
      P[ 246] <= 9'b110000000; // Load the target box with 0
      P[ 247] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 248] <= 9'b000000000; // Load the constant box with 0
      P[ 249] <= 9'b101000001; // Load the source box with 1
      P[ 250] <= 9'b110000110; // Load the target box with 6
      P[ 251] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 252] <= 9'b000001001; // Load the constant box with 9
      P[ 253] <= 9'b101000110; // Load the source box with 6
      P[ 254] <= 9'b110000000; // Load the target box with 0
      P[ 255] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 256] <= 9'b000001111; // Load the constant box with 15
      P[ 257] <= 9'b101000110; // Load the source box with 6
      P[ 258] <= 9'b110000000; // Load the target box with 0
      P[ 259] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 260] <= 9'b000000000; // Load the constant box with 0
      P[ 261] <= 9'b101000001; // Load the source box with 1
      P[ 262] <= 9'b110000111; // Load the target box with 7
      P[ 263] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 264] <= 9'b000001010; // Load the constant box with 10
      P[ 265] <= 9'b101000111; // Load the source box with 7
      P[ 266] <= 9'b110000000; // Load the target box with 0
      P[ 267] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 268] <= 9'b000001111; // Load the constant box with 15
      P[ 269] <= 9'b101000111; // Load the source box with 7
      P[ 270] <= 9'b110000000; // Load the target box with 0
      P[ 271] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 272] <= 9'b000000000; // Load the constant box with 0
      P[ 273] <= 9'b101000001; // Load the source box with 1
      P[ 274] <= 9'b110001000; // Load the target box with 8
      P[ 275] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 276] <= 9'b000001011; // Load the constant box with 11
      P[ 277] <= 9'b101001000; // Load the source box with 8
      P[ 278] <= 9'b110000000; // Load the target box with 0
      P[ 279] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 280] <= 9'b000001111; // Load the constant box with 15
      P[ 281] <= 9'b101001000; // Load the source box with 8
      P[ 282] <= 9'b110000000; // Load the target box with 0
      P[ 283] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 284] <= 9'b000000000; // Load the constant box with 0
      P[ 285] <= 9'b101000001; // Load the source box with 1
      P[ 286] <= 9'b110001001; // Load the target box with 9
      P[ 287] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 288] <= 9'b000001100; // Load the constant box with 12
      P[ 289] <= 9'b101001001; // Load the source box with 9
      P[ 290] <= 9'b110000000; // Load the target box with 0
      P[ 291] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 292] <= 9'b000001111; // Load the constant box with 15
      P[ 293] <= 9'b101001001; // Load the source box with 9
      P[ 294] <= 9'b110000000; // Load the target box with 0
      P[ 295] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 296] <= 9'b000000000; // Load the constant box with 0
      P[ 297] <= 9'b101000001; // Load the source box with 1
      P[ 298] <= 9'b110001010; // Load the target box with 10
      P[ 299] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 300] <= 9'b000001101; // Load the constant box with 13
      P[ 301] <= 9'b101001010; // Load the source box with 10
      P[ 302] <= 9'b110000000; // Load the target box with 0
      P[ 303] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 304] <= 9'b000001111; // Load the constant box with 15
      P[ 305] <= 9'b101001010; // Load the source box with 10
      P[ 306] <= 9'b110000000; // Load the target box with 0
      P[ 307] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 308] <= 9'b000000000; // Load the constant box with 0
      P[ 309] <= 9'b101000001; // Load the source box with 1
      P[ 310] <= 9'b110001011; // Load the target box with 11
      P[ 311] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 312] <= 9'b000001110; // Load the constant box with 14
      P[ 313] <= 9'b101001011; // Load the source box with 11
      P[ 314] <= 9'b110000000; // Load the target box with 0
      P[ 315] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 316] <= 9'b000001111; // Load the constant box with 15
      P[ 317] <= 9'b101001011; // Load the source box with 11
      P[ 318] <= 9'b110000000; // Load the target box with 0
      P[ 319] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 320] <= 9'b000000000; // Load the constant box with 0
      P[ 321] <= 9'b101000001; // Load the source box with 1
      P[ 322] <= 9'b110001100; // Load the target box with 12
      P[ 323] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 324] <= 9'b000001111; // Load the constant box with 15
      P[ 325] <= 9'b101001100; // Load the source box with 12
      P[ 326] <= 9'b110000000; // Load the target box with 0
      P[ 327] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 328] <= 9'b000001111; // Load the constant box with 15
      P[ 329] <= 9'b101001100; // Load the source box with 12
      P[ 330] <= 9'b110000000; // Load the target box with 0
      P[ 331] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 332] <= 9'b000000000; // Load the constant box with 0
      P[ 333] <= 9'b101000001; // Load the source box with 1
      P[ 334] <= 9'b110001101; // Load the target box with 13
      P[ 335] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 336] <= 9'b000000101; // Load the constant box with 5
      P[ 337] <= 9'b101001101; // Load the source box with 13
      P[ 338] <= 9'b110000000; // Load the target box with 0
      P[ 339] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 340] <= 9'b000001001; // Load the constant box with 9
      P[ 341] <= 9'b101001101; // Load the source box with 13
      P[ 342] <= 9'b110000000; // Load the target box with 0
      P[ 343] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 344] <= 9'b000000001; // Load the constant box with 1
      P[ 345] <= 9'b101001101; // Load the source box with 13
      P[ 346] <= 9'b110000000; // Load the target box with 0
      P[ 347] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 348] <= 9'b000000000; // Load the constant box with 0
      P[ 349] <= 9'b101000001; // Load the source box with 1
      P[ 350] <= 9'b110001110; // Load the target box with 14
      P[ 351] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 352] <= 9'b000001000; // Load the constant box with 8
      P[ 353] <= 9'b101001110; // Load the source box with 14
      P[ 354] <= 9'b110000000; // Load the target box with 0
      P[ 355] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 356] <= 9'b000001101; // Load the constant box with 13
      P[ 357] <= 9'b101001110; // Load the source box with 14
      P[ 358] <= 9'b110000000; // Load the target box with 0
      P[ 359] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 360] <= 9'b000000101; // Load the constant box with 5
      P[ 361] <= 9'b101001110; // Load the source box with 14
      P[ 362] <= 9'b110000000; // Load the target box with 0
      P[ 363] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 364] <= 9'b000000000; // Load the constant box with 0
      P[ 365] <= 9'b101000001; // Load the source box with 1
      P[ 366] <= 9'b110001111; // Load the target box with 15
      P[ 367] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 368] <= 9'b000001111; // Load the constant box with 15
      P[ 369] <= 9'b101001111; // Load the source box with 15
      P[ 370] <= 9'b110000000; // Load the target box with 0
      P[ 371] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 372] <= 9'b000001100; // Load the constant box with 12
      P[ 373] <= 9'b101001111; // Load the source box with 15
      P[ 374] <= 9'b110000000; // Load the target box with 0
      P[ 375] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 376] <= 9'b000000000; // Load the constant box with 0
      P[ 377] <= 9'b101001111; // Load the source box with 15
      P[ 378] <= 9'b110001110; // Load the target box with 14
      P[ 379] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 380] <= 9'b000000000; // Load the constant box with 0
      P[ 381] <= 9'b101000010; // Load the source box with 2
      P[ 382] <= 9'b110001111; // Load the target box with 15
      P[ 383] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 384] <= 9'b000000000; // Load the constant box with 0
      P[ 385] <= 9'b101000011; // Load the source box with 3
      P[ 386] <= 9'b110001111; // Load the target box with 15
      P[ 387] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 388] <= 9'b000000000; // Load the constant box with 0
      P[ 389] <= 9'b101000100; // Load the source box with 4
      P[ 390] <= 9'b110001111; // Load the target box with 15
      P[ 391] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 392] <= 9'b000000000; // Load the constant box with 0
      P[ 393] <= 9'b101000101; // Load the source box with 5
      P[ 394] <= 9'b110001111; // Load the target box with 15
      P[ 395] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 396] <= 9'b000000000; // Load the constant box with 0
      P[ 397] <= 9'b101000110; // Load the source box with 6
      P[ 398] <= 9'b110001111; // Load the target box with 15
      P[ 399] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 400] <= 9'b000000000; // Load the constant box with 0
      P[ 401] <= 9'b101000111; // Load the source box with 7
      P[ 402] <= 9'b110001111; // Load the target box with 15
      P[ 403] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 404] <= 9'b000000000; // Load the constant box with 0
      P[ 405] <= 9'b101001000; // Load the source box with 8
      P[ 406] <= 9'b110001111; // Load the target box with 15
      P[ 407] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 408] <= 9'b000000001; // Load the constant box with 1
      P[ 409] <= 9'b101000000; // Load the source box with 0
      P[ 410] <= 9'b110000000; // Load the target box with 0
      P[ 411] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 412] <= 9'b000000000; // Load the constant box with 0
      P[ 413] <= 9'b101001111; // Load the source box with 15
      P[ 414] <= 9'b110000000; // Load the target box with 0
      P[ 415] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 416] <= 9'b011110111; // Load the constant box with 247
      P[ 417] <= 9'b101000000; // Load the source box with 0
      P[ 418] <= 9'b110000000; // Load the target box with 0
      P[ 419] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 420] <= 9'b000000000; // Load the constant box with 0
      P[ 421] <= 9'b101000000; // Load the source box with 0
      P[ 422] <= 9'b110000001; // Load the target box with 1
      P[ 423] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 424] <= 9'b000000000; // Load the constant box with 0
      P[ 425] <= 9'b101000000; // Load the source box with 0
      P[ 426] <= 9'b110001101; // Load the target box with 13
      P[ 427] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 428] <= 9'b000000000; // Load the constant box with 0
      P[ 429] <= 9'b101000010; // Load the source box with 2
      P[ 430] <= 9'b110001111; // Load the target box with 15
      P[ 431] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 432] <= 9'b000000000; // Load the constant box with 0
      P[ 433] <= 9'b101000011; // Load the source box with 3
      P[ 434] <= 9'b110001111; // Load the target box with 15
      P[ 435] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 436] <= 9'b000000000; // Load the constant box with 0
      P[ 437] <= 9'b101000100; // Load the source box with 4
      P[ 438] <= 9'b110001111; // Load the target box with 15
      P[ 439] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 440] <= 9'b000000000; // Load the constant box with 0
      P[ 441] <= 9'b101000101; // Load the source box with 5
      P[ 442] <= 9'b110001111; // Load the target box with 15
      P[ 443] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 444] <= 9'b000000000; // Load the constant box with 0
      P[ 445] <= 9'b101001001; // Load the source box with 9
      P[ 446] <= 9'b110001111; // Load the target box with 15
      P[ 447] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 448] <= 9'b000000000; // Load the constant box with 0
      P[ 449] <= 9'b101001010; // Load the source box with 10
      P[ 450] <= 9'b110001111; // Load the target box with 15
      P[ 451] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 452] <= 9'b000000000; // Load the constant box with 0
      P[ 453] <= 9'b101001011; // Load the source box with 11
      P[ 454] <= 9'b110001111; // Load the target box with 15
      P[ 455] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 456] <= 9'b000000001; // Load the constant box with 1
      P[ 457] <= 9'b101000000; // Load the source box with 0
      P[ 458] <= 9'b110000000; // Load the target box with 0
      P[ 459] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 460] <= 9'b000000000; // Load the constant box with 0
      P[ 461] <= 9'b101001111; // Load the source box with 15
      P[ 462] <= 9'b110000000; // Load the target box with 0
      P[ 463] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 464] <= 9'b011111000; // Load the constant box with 248
      P[ 465] <= 9'b101000000; // Load the source box with 0
      P[ 466] <= 9'b110000000; // Load the target box with 0
      P[ 467] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 468] <= 9'b000000000; // Load the constant box with 0
      P[ 469] <= 9'b101000000; // Load the source box with 0
      P[ 470] <= 9'b110000001; // Load the target box with 1
      P[ 471] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 472] <= 9'b000000100; // Load the constant box with 4
      P[ 473] <= 9'b101000000; // Load the source box with 0
      P[ 474] <= 9'b110000000; // Load the target box with 0
      P[ 475] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 476] <= 9'b000000000; // Load the constant box with 0
      P[ 477] <= 9'b101000000; // Load the source box with 0
      P[ 478] <= 9'b110001110; // Load the target box with 14
      P[ 479] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 480] <= 9'b000000000; // Load the constant box with 0
      P[ 481] <= 9'b101000010; // Load the source box with 2
      P[ 482] <= 9'b110001111; // Load the target box with 15
      P[ 483] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 484] <= 9'b000000000; // Load the constant box with 0
      P[ 485] <= 9'b101000011; // Load the source box with 3
      P[ 486] <= 9'b110001111; // Load the target box with 15
      P[ 487] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 488] <= 9'b000000000; // Load the constant box with 0
      P[ 489] <= 9'b101000110; // Load the source box with 6
      P[ 490] <= 9'b110001111; // Load the target box with 15
      P[ 491] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 492] <= 9'b000000000; // Load the constant box with 0
      P[ 493] <= 9'b101000111; // Load the source box with 7
      P[ 494] <= 9'b110001111; // Load the target box with 15
      P[ 495] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 496] <= 9'b000000000; // Load the constant box with 0
      P[ 497] <= 9'b101001001; // Load the source box with 9
      P[ 498] <= 9'b110001111; // Load the target box with 15
      P[ 499] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 500] <= 9'b000000000; // Load the constant box with 0
      P[ 501] <= 9'b101001010; // Load the source box with 10
      P[ 502] <= 9'b110001111; // Load the target box with 15
      P[ 503] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 504] <= 9'b000000000; // Load the constant box with 0
      P[ 505] <= 9'b101001100; // Load the source box with 12
      P[ 506] <= 9'b110001111; // Load the target box with 15
      P[ 507] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 508] <= 9'b000000001; // Load the constant box with 1
      P[ 509] <= 9'b101000000; // Load the source box with 0
      P[ 510] <= 9'b110000000; // Load the target box with 0
      P[ 511] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 512] <= 9'b000000000; // Load the constant box with 0
      P[ 513] <= 9'b101001111; // Load the source box with 15
      P[ 514] <= 9'b110000000; // Load the target box with 0
      P[ 515] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 516] <= 9'b011111001; // Load the constant box with 249
      P[ 517] <= 9'b101000000; // Load the source box with 0
      P[ 518] <= 9'b110000000; // Load the target box with 0
      P[ 519] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 520] <= 9'b000000000; // Load the constant box with 0
      P[ 521] <= 9'b101000000; // Load the source box with 0
      P[ 522] <= 9'b110000001; // Load the target box with 1
      P[ 523] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 524] <= 9'b000000010; // Load the constant box with 2
      P[ 525] <= 9'b101000000; // Load the source box with 0
      P[ 526] <= 9'b110000000; // Load the target box with 0
      P[ 527] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 528] <= 9'b000000000; // Load the constant box with 0
      P[ 529] <= 9'b101000000; // Load the source box with 0
      P[ 530] <= 9'b110001110; // Load the target box with 14
      P[ 531] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 532] <= 9'b000000000; // Load the constant box with 0
      P[ 533] <= 9'b101000010; // Load the source box with 2
      P[ 534] <= 9'b110001111; // Load the target box with 15
      P[ 535] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 536] <= 9'b000000000; // Load the constant box with 0
      P[ 537] <= 9'b101000100; // Load the source box with 4
      P[ 538] <= 9'b110001111; // Load the target box with 15
      P[ 539] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 540] <= 9'b000000000; // Load the constant box with 0
      P[ 541] <= 9'b101000110; // Load the source box with 6
      P[ 542] <= 9'b110001111; // Load the target box with 15
      P[ 543] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 544] <= 9'b000000000; // Load the constant box with 0
      P[ 545] <= 9'b101001000; // Load the source box with 8
      P[ 546] <= 9'b110001111; // Load the target box with 15
      P[ 547] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 548] <= 9'b000000000; // Load the constant box with 0
      P[ 549] <= 9'b101001001; // Load the source box with 9
      P[ 550] <= 9'b110001111; // Load the target box with 15
      P[ 551] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 552] <= 9'b000000000; // Load the constant box with 0
      P[ 553] <= 9'b101001011; // Load the source box with 11
      P[ 554] <= 9'b110001111; // Load the target box with 15
      P[ 555] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 556] <= 9'b000000000; // Load the constant box with 0
      P[ 557] <= 9'b101001100; // Load the source box with 12
      P[ 558] <= 9'b110001111; // Load the target box with 15
      P[ 559] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 560] <= 9'b000000001; // Load the constant box with 1
      P[ 561] <= 9'b101000000; // Load the source box with 0
      P[ 562] <= 9'b110000000; // Load the target box with 0
      P[ 563] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 564] <= 9'b000000000; // Load the constant box with 0
      P[ 565] <= 9'b101001111; // Load the source box with 15
      P[ 566] <= 9'b110000000; // Load the target box with 0
      P[ 567] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 568] <= 9'b011111010; // Load the constant box with 250
      P[ 569] <= 9'b101000000; // Load the source box with 0
      P[ 570] <= 9'b110000000; // Load the target box with 0
      P[ 571] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 572] <= 9'b000000000; // Load the constant box with 0
      P[ 573] <= 9'b101000000; // Load the source box with 0
      P[ 574] <= 9'b110000001; // Load the target box with 1
      P[ 575] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 576] <= 9'b000000001; // Load the constant box with 1
      P[ 577] <= 9'b101000000; // Load the source box with 0
      P[ 578] <= 9'b110000000; // Load the target box with 0
      P[ 579] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 580] <= 9'b000000000; // Load the constant box with 0
      P[ 581] <= 9'b101000000; // Load the source box with 0
      P[ 582] <= 9'b110001110; // Load the target box with 14
      P[ 583] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 584] <= 9'b000000000; // Load the constant box with 0
      P[ 585] <= 9'b101000010; // Load the source box with 2
      P[ 586] <= 9'b110000001; // Load the target box with 1
      P[ 587] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 588] <= 9'b000000000; // Load the constant box with 0
      P[ 589] <= 9'b101000011; // Load the source box with 3
      P[ 590] <= 9'b110000001; // Load the target box with 1
      P[ 591] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 592] <= 9'b000000000; // Load the constant box with 0
      P[ 593] <= 9'b101000100; // Load the source box with 4
      P[ 594] <= 9'b110000001; // Load the target box with 1
      P[ 595] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 596] <= 9'b000000000; // Load the constant box with 0
      P[ 597] <= 9'b101000101; // Load the source box with 5
      P[ 598] <= 9'b110000001; // Load the target box with 1
      P[ 599] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 600] <= 9'b000000000; // Load the constant box with 0
      P[ 601] <= 9'b101000110; // Load the source box with 6
      P[ 602] <= 9'b110000001; // Load the target box with 1
      P[ 603] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 604] <= 9'b000000000; // Load the constant box with 0
      P[ 605] <= 9'b101000111; // Load the source box with 7
      P[ 606] <= 9'b110000001; // Load the target box with 1
      P[ 607] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 608] <= 9'b000000000; // Load the constant box with 0
      P[ 609] <= 9'b101001000; // Load the source box with 8
      P[ 610] <= 9'b110000001; // Load the target box with 1
      P[ 611] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 612] <= 9'b000000000; // Load the constant box with 0
      P[ 613] <= 9'b101001001; // Load the source box with 9
      P[ 614] <= 9'b110000001; // Load the target box with 1
      P[ 615] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 616] <= 9'b000000000; // Load the constant box with 0
      P[ 617] <= 9'b101001010; // Load the source box with 10
      P[ 618] <= 9'b110000001; // Load the target box with 1
      P[ 619] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 620] <= 9'b000000000; // Load the constant box with 0
      P[ 621] <= 9'b101001011; // Load the source box with 11
      P[ 622] <= 9'b110000001; // Load the target box with 1
      P[ 623] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 624] <= 9'b000000000; // Load the constant box with 0
      P[ 625] <= 9'b101001100; // Load the source box with 12
      P[ 626] <= 9'b110000001; // Load the target box with 1
      P[ 627] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 628] <= 9'b000000001; // Load the constant box with 1
      P[ 629] <= 9'b101000000; // Load the source box with 0
      P[ 630] <= 9'b110000000; // Load the target box with 0
      P[ 631] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 632] <= 9'b000000000; // Load the constant box with 0
      P[ 633] <= 9'b101000001; // Load the source box with 1
      P[ 634] <= 9'b110000000; // Load the target box with 0
      P[ 635] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 636] <= 9'b011110110; // Load the constant box with 246
      P[ 637] <= 9'b101000000; // Load the source box with 0
      P[ 638] <= 9'b110000000; // Load the target box with 0
      P[ 639] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 640] <= 9'b000000000; // Load the constant box with 0
      P[ 641] <= 9'b101000000; // Load the source box with 0
      P[ 642] <= 9'b110001110; // Load the target box with 14
      P[ 643] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 644] <= 9'b011111100; // Load the constant box with 252
      P[ 645] <= 9'b101001101; // Load the source box with 13
      P[ 646] <= 9'b110000000; // Load the target box with 0
      P[ 647] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 648] <= 9'b011111011; // Load the constant box with 251
      P[ 649] <= 9'b101001110; // Load the source box with 14
      P[ 650] <= 9'b110000000; // Load the target box with 0
      P[ 651] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 652] <= 9'b000000000; // Load the constant box with 0
      P[ 653] <= 9'b101000000; // Load the source box with 0
      P[ 654] <= 9'b110000000; // Load the target box with 0
      P[ 655] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 656] <= 9'b011110110; // Load the constant box with 246
      P[ 657] <= 9'b101000001; // Load the source box with 1
      P[ 658] <= 9'b110000000; // Load the target box with 0
      P[ 659] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 660] <= 9'b011110001; // Load the constant box with 241
      P[ 661] <= 9'b101000010; // Load the source box with 2
      P[ 662] <= 9'b110000000; // Load the target box with 0
      P[ 663] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 664] <= 9'b000000000; // Load the constant box with 0
      P[ 665] <= 9'b101000010; // Load the source box with 2
      P[ 666] <= 9'b110000001; // Load the target box with 1
      P[ 667] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 668] <= 9'b000000100; // Load the constant box with 4
      P[ 669] <= 9'b101000001; // Load the source box with 1
      P[ 670] <= 9'b110000000; // Load the target box with 0
      P[ 671] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 672] <= 9'b000000000; // Load the constant box with 0
      P[ 673] <= 9'b101000001; // Load the source box with 1
      P[ 674] <= 9'b110000000; // Load the target box with 0
      P[ 675] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 676] <= 9'b011110111; // Load the constant box with 247
      P[ 677] <= 9'b101000001; // Load the source box with 1
      P[ 678] <= 9'b110000000; // Load the target box with 0
      P[ 679] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 680] <= 9'b011110010; // Load the constant box with 242
      P[ 681] <= 9'b101000010; // Load the source box with 2
      P[ 682] <= 9'b110000000; // Load the target box with 0
      P[ 683] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 684] <= 9'b000000000; // Load the constant box with 0
      P[ 685] <= 9'b101000010; // Load the source box with 2
      P[ 686] <= 9'b110000001; // Load the target box with 1
      P[ 687] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 688] <= 9'b000000011; // Load the constant box with 3
      P[ 689] <= 9'b101000001; // Load the source box with 1
      P[ 690] <= 9'b110000000; // Load the target box with 0
      P[ 691] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 692] <= 9'b000000000; // Load the constant box with 0
      P[ 693] <= 9'b101000001; // Load the source box with 1
      P[ 694] <= 9'b110000000; // Load the target box with 0
      P[ 695] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 696] <= 9'b011111000; // Load the constant box with 248
      P[ 697] <= 9'b101000001; // Load the source box with 1
      P[ 698] <= 9'b110000000; // Load the target box with 0
      P[ 699] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 700] <= 9'b011110011; // Load the constant box with 243
      P[ 701] <= 9'b101000010; // Load the source box with 2
      P[ 702] <= 9'b110000000; // Load the target box with 0
      P[ 703] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 704] <= 9'b000000000; // Load the constant box with 0
      P[ 705] <= 9'b101000010; // Load the source box with 2
      P[ 706] <= 9'b110000001; // Load the target box with 1
      P[ 707] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 708] <= 9'b000000010; // Load the constant box with 2
      P[ 709] <= 9'b101000001; // Load the source box with 1
      P[ 710] <= 9'b110000000; // Load the target box with 0
      P[ 711] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 712] <= 9'b000000000; // Load the constant box with 0
      P[ 713] <= 9'b101000001; // Load the source box with 1
      P[ 714] <= 9'b110000000; // Load the target box with 0
      P[ 715] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 716] <= 9'b011111001; // Load the constant box with 249
      P[ 717] <= 9'b101000001; // Load the source box with 1
      P[ 718] <= 9'b110000000; // Load the target box with 0
      P[ 719] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 720] <= 9'b011110100; // Load the constant box with 244
      P[ 721] <= 9'b101000010; // Load the source box with 2
      P[ 722] <= 9'b110000000; // Load the target box with 0
      P[ 723] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 724] <= 9'b000000000; // Load the constant box with 0
      P[ 725] <= 9'b101000010; // Load the source box with 2
      P[ 726] <= 9'b110000001; // Load the target box with 1
      P[ 727] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 728] <= 9'b000000001; // Load the constant box with 1
      P[ 729] <= 9'b101000001; // Load the source box with 1
      P[ 730] <= 9'b110000000; // Load the target box with 0
      P[ 731] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 732] <= 9'b000000000; // Load the constant box with 0
      P[ 733] <= 9'b101000001; // Load the source box with 1
      P[ 734] <= 9'b110000000; // Load the target box with 0
      P[ 735] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 736] <= 9'b011111010; // Load the constant box with 250
      P[ 737] <= 9'b101000001; // Load the source box with 1
      P[ 738] <= 9'b110000000; // Load the target box with 0
      P[ 739] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 740] <= 9'b011110101; // Load the constant box with 245
      P[ 741] <= 9'b101000010; // Load the source box with 2
      P[ 742] <= 9'b110000000; // Load the target box with 0
      P[ 743] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 744] <= 9'b000000000; // Load the constant box with 0
      P[ 745] <= 9'b101000010; // Load the source box with 2
      P[ 746] <= 9'b110000001; // Load the target box with 1
      P[ 747] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 748] <= 9'b000000000; // Load the constant box with 0
      P[ 749] <= 9'b101000001; // Load the source box with 1
      P[ 750] <= 9'b110000000; // Load the target box with 0
      P[ 751] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 752] <= 9'b000000000; // Load the constant box with 0
      P[ 753] <= 9'b101000000; // Load the source box with 0
      P[ 754] <= 9'b110000000; // Load the target box with 0
      P[ 755] <= 9'b111001110; // not: Invert the bits in a register
      P[ 756] <= 9'b000011111; // Load the constant box with 31
      P[ 757] <= 9'b101000001; // Load the source box with 1
      P[ 758] <= 9'b110000000; // Load the target box with 0
      P[ 759] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 760] <= 9'b000000000; // Load the constant box with 0
      P[ 761] <= 9'b101000001; // Load the source box with 1
      P[ 762] <= 9'b110000000; // Load the target box with 0
      P[ 763] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 764] <= 9'b010010010; // Load the constant box with 146
      P[ 765] <= 9'b101000000; // Load the source box with 0
      P[ 766] <= 9'b110000000; // Load the target box with 0
      P[ 767] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 768] <= 9'b000000000; // Load the constant box with 0
      P[ 769] <= 9'b101000000; // Load the source box with 0
      P[ 770] <= 9'b110000001; // Load the target box with 1
      P[ 771] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 772] <= 9'b000011111; // Load the constant box with 31
      P[ 773] <= 9'b101000010; // Load the source box with 2
      P[ 774] <= 9'b110000000; // Load the target box with 0
      P[ 775] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 776] <= 9'b000000000; // Load the constant box with 0
      P[ 777] <= 9'b101000010; // Load the source box with 2
      P[ 778] <= 9'b110000001; // Load the target box with 1
      P[ 779] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 780] <= 9'b000001101; // Load the constant box with 13
      P[ 781] <= 9'b101000000; // Load the source box with 0
      P[ 782] <= 9'b110000000; // Load the target box with 0
      P[ 783] <= 9'b111001001; // label: Create and set a label
      P[ 784] <= 9'b001100100; // Load the constant box with 100
      P[ 785] <= 9'b101000001; // Load the source box with 1
      P[ 786] <= 9'b110000000; // Load the target box with 0
      P[ 787] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 788] <= 9'b011111110; // Load the constant box with 254
      P[ 789] <= 9'b101000011; // Load the source box with 3
      P[ 790] <= 9'b110000000; // Load the target box with 0
      P[ 791] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 792] <= 9'b000000100; // Load the constant box with 4
      P[ 793] <= 9'b101000011; // Load the source box with 3
      P[ 794] <= 9'b110000000; // Load the target box with 0
      P[ 795] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[ 796] <= 9'b011111110; // Load the constant box with 254
      P[ 797] <= 9'b101000011; // Load the source box with 3
      P[ 798] <= 9'b110000000; // Load the target box with 0
      P[ 799] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 800] <= 9'b000000011; // Load the constant box with 3
      P[ 801] <= 9'b101000000; // Load the source box with 0
      P[ 802] <= 9'b110000000; // Load the target box with 0
      P[ 803] <= 9'b111001001; // label: Set a label
      P[ 804] <= 9'b000000000; // Load the constant box with 0
      P[ 805] <= 9'b101000000; // Load the source box with 0
      P[ 806] <= 9'b110000001; // Load the target box with 1
      P[ 807] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 808] <= 9'b000001110; // Load the constant box with 14
      P[ 809] <= 9'b101000010; // Load the source box with 2
      P[ 810] <= 9'b110000000; // Load the target box with 0
      P[ 811] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 812] <= 9'b000000000; // Load the constant box with 0
      P[ 813] <= 9'b101000010; // Load the source box with 2
      P[ 814] <= 9'b110000001; // Load the target box with 1
      P[ 815] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 816] <= 9'b000001101; // Load the constant box with 13
      P[ 817] <= 9'b101000000; // Load the source box with 0
      P[ 818] <= 9'b110000000; // Load the target box with 0
      P[ 819] <= 9'b111001001; // label: Create and set a label
      P[ 820] <= 9'b001101001; // Load the constant box with 105
      P[ 821] <= 9'b101000001; // Load the source box with 1
      P[ 822] <= 9'b110000000; // Load the target box with 0
      P[ 823] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 824] <= 9'b011111110; // Load the constant box with 254
      P[ 825] <= 9'b101000011; // Load the source box with 3
      P[ 826] <= 9'b110000000; // Load the target box with 0
      P[ 827] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 828] <= 9'b000000010; // Load the constant box with 2
      P[ 829] <= 9'b101000011; // Load the source box with 3
      P[ 830] <= 9'b110000000; // Load the target box with 0
      P[ 831] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[ 832] <= 9'b011111110; // Load the constant box with 254
      P[ 833] <= 9'b101000011; // Load the source box with 3
      P[ 834] <= 9'b110000000; // Load the target box with 0
      P[ 835] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 836] <= 9'b000000100; // Load the constant box with 4
      P[ 837] <= 9'b101000000; // Load the source box with 0
      P[ 838] <= 9'b110000000; // Load the target box with 0
      P[ 839] <= 9'b111001001; // label: Set a label
      P[ 840] <= 9'b000000000; // Load the constant box with 0
      P[ 841] <= 9'b101000000; // Load the source box with 0
      P[ 842] <= 9'b110000001; // Load the target box with 1
      P[ 843] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 844] <= 9'b000001101; // Load the constant box with 13
      P[ 845] <= 9'b101000010; // Load the source box with 2
      P[ 846] <= 9'b110000000; // Load the target box with 0
      P[ 847] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 848] <= 9'b000000000; // Load the constant box with 0
      P[ 849] <= 9'b101000010; // Load the source box with 2
      P[ 850] <= 9'b110000001; // Load the target box with 1
      P[ 851] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 852] <= 9'b000001101; // Load the constant box with 13
      P[ 853] <= 9'b101000000; // Load the source box with 0
      P[ 854] <= 9'b110000000; // Load the target box with 0
      P[ 855] <= 9'b111001001; // label: Create and set a label
      P[ 856] <= 9'b001101101; // Load the constant box with 109
      P[ 857] <= 9'b101000001; // Load the source box with 1
      P[ 858] <= 9'b110000000; // Load the target box with 0
      P[ 859] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 860] <= 9'b011111110; // Load the constant box with 254
      P[ 861] <= 9'b101000011; // Load the source box with 3
      P[ 862] <= 9'b110000000; // Load the target box with 0
      P[ 863] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 864] <= 9'b000000001; // Load the constant box with 1
      P[ 865] <= 9'b101000011; // Load the source box with 3
      P[ 866] <= 9'b110000000; // Load the target box with 0
      P[ 867] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[ 868] <= 9'b011111110; // Load the constant box with 254
      P[ 869] <= 9'b101000011; // Load the source box with 3
      P[ 870] <= 9'b110000000; // Load the target box with 0
      P[ 871] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 872] <= 9'b000000101; // Load the constant box with 5
      P[ 873] <= 9'b101000000; // Load the source box with 0
      P[ 874] <= 9'b110000000; // Load the target box with 0
      P[ 875] <= 9'b111001001; // label: Set a label
      P[ 876] <= 9'b000000000; // Load the constant box with 0
      P[ 877] <= 9'b101000000; // Load the source box with 0
      P[ 878] <= 9'b110000001; // Load the target box with 1
      P[ 879] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 880] <= 9'b000011100; // Load the constant box with 28
      P[ 881] <= 9'b101000010; // Load the source box with 2
      P[ 882] <= 9'b110000000; // Load the target box with 0
      P[ 883] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 884] <= 9'b000000000; // Load the constant box with 0
      P[ 885] <= 9'b101000010; // Load the source box with 2
      P[ 886] <= 9'b110000001; // Load the target box with 1
      P[ 887] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 888] <= 9'b000001101; // Load the constant box with 13
      P[ 889] <= 9'b101000000; // Load the source box with 0
      P[ 890] <= 9'b110000000; // Load the target box with 0
      P[ 891] <= 9'b111001001; // label: Create and set a label
      P[ 892] <= 9'b001110010; // Load the constant box with 114
      P[ 893] <= 9'b101000001; // Load the source box with 1
      P[ 894] <= 9'b110000000; // Load the target box with 0
      P[ 895] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 896] <= 9'b011111101; // Load the constant box with 253
      P[ 897] <= 9'b101000011; // Load the source box with 3
      P[ 898] <= 9'b110000000; // Load the target box with 0
      P[ 899] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 900] <= 9'b010000000; // Load the constant box with 128
      P[ 901] <= 9'b101000011; // Load the source box with 3
      P[ 902] <= 9'b110000000; // Load the target box with 0
      P[ 903] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[ 904] <= 9'b011111101; // Load the constant box with 253
      P[ 905] <= 9'b101000011; // Load the source box with 3
      P[ 906] <= 9'b110000000; // Load the target box with 0
      P[ 907] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 908] <= 9'b000000110; // Load the constant box with 6
      P[ 909] <= 9'b101000000; // Load the source box with 0
      P[ 910] <= 9'b110000000; // Load the target box with 0
      P[ 911] <= 9'b111001001; // label: Set a label
      P[ 912] <= 9'b000000000; // Load the constant box with 0
      P[ 913] <= 9'b101000000; // Load the source box with 0
      P[ 914] <= 9'b110000001; // Load the target box with 1
      P[ 915] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 916] <= 9'b000001011; // Load the constant box with 11
      P[ 917] <= 9'b101000010; // Load the source box with 2
      P[ 918] <= 9'b110000000; // Load the target box with 0
      P[ 919] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 920] <= 9'b000000000; // Load the constant box with 0
      P[ 921] <= 9'b101000010; // Load the source box with 2
      P[ 922] <= 9'b110000001; // Load the target box with 1
      P[ 923] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 924] <= 9'b000001101; // Load the constant box with 13
      P[ 925] <= 9'b101000000; // Load the source box with 0
      P[ 926] <= 9'b110000000; // Load the target box with 0
      P[ 927] <= 9'b111001001; // label: Create and set a label
      P[ 928] <= 9'b001110110; // Load the constant box with 118
      P[ 929] <= 9'b101000001; // Load the source box with 1
      P[ 930] <= 9'b110000000; // Load the target box with 0
      P[ 931] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 932] <= 9'b011111101; // Load the constant box with 253
      P[ 933] <= 9'b101000011; // Load the source box with 3
      P[ 934] <= 9'b110000000; // Load the target box with 0
      P[ 935] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 936] <= 9'b001000000; // Load the constant box with 64
      P[ 937] <= 9'b101000011; // Load the source box with 3
      P[ 938] <= 9'b110000000; // Load the target box with 0
      P[ 939] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[ 940] <= 9'b011111101; // Load the constant box with 253
      P[ 941] <= 9'b101000011; // Load the source box with 3
      P[ 942] <= 9'b110000000; // Load the target box with 0
      P[ 943] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 944] <= 9'b000000111; // Load the constant box with 7
      P[ 945] <= 9'b101000000; // Load the source box with 0
      P[ 946] <= 9'b110000000; // Load the target box with 0
      P[ 947] <= 9'b111001001; // label: Set a label
      P[ 948] <= 9'b000000000; // Load the constant box with 0
      P[ 949] <= 9'b101000000; // Load the source box with 0
      P[ 950] <= 9'b110000001; // Load the target box with 1
      P[ 951] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 952] <= 9'b000011010; // Load the constant box with 26
      P[ 953] <= 9'b101000010; // Load the source box with 2
      P[ 954] <= 9'b110000000; // Load the target box with 0
      P[ 955] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 956] <= 9'b000000000; // Load the constant box with 0
      P[ 957] <= 9'b101000010; // Load the source box with 2
      P[ 958] <= 9'b110000001; // Load the target box with 1
      P[ 959] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 960] <= 9'b000001101; // Load the constant box with 13
      P[ 961] <= 9'b101000000; // Load the source box with 0
      P[ 962] <= 9'b110000000; // Load the target box with 0
      P[ 963] <= 9'b111001001; // label: Create and set a label
      P[ 964] <= 9'b001111011; // Load the constant box with 123
      P[ 965] <= 9'b101000001; // Load the source box with 1
      P[ 966] <= 9'b110000000; // Load the target box with 0
      P[ 967] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 968] <= 9'b011111101; // Load the constant box with 253
      P[ 969] <= 9'b101000011; // Load the source box with 3
      P[ 970] <= 9'b110000000; // Load the target box with 0
      P[ 971] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[ 972] <= 9'b000100000; // Load the constant box with 32
      P[ 973] <= 9'b101000011; // Load the source box with 3
      P[ 974] <= 9'b110000000; // Load the target box with 0
      P[ 975] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[ 976] <= 9'b011111101; // Load the constant box with 253
      P[ 977] <= 9'b101000011; // Load the source box with 3
      P[ 978] <= 9'b110000000; // Load the target box with 0
      P[ 979] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 980] <= 9'b000001000; // Load the constant box with 8
      P[ 981] <= 9'b101000000; // Load the source box with 0
      P[ 982] <= 9'b110000000; // Load the target box with 0
      P[ 983] <= 9'b111001001; // label: Set a label
      P[ 984] <= 9'b000000000; // Load the constant box with 0
      P[ 985] <= 9'b101000000; // Load the source box with 0
      P[ 986] <= 9'b110000001; // Load the target box with 1
      P[ 987] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 988] <= 9'b000011001; // Load the constant box with 25
      P[ 989] <= 9'b101000010; // Load the source box with 2
      P[ 990] <= 9'b110000000; // Load the target box with 0
      P[ 991] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 992] <= 9'b000000000; // Load the constant box with 0
      P[ 993] <= 9'b101000010; // Load the source box with 2
      P[ 994] <= 9'b110000001; // Load the target box with 1
      P[ 995] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 996] <= 9'b000001101; // Load the constant box with 13
      P[ 997] <= 9'b101000000; // Load the source box with 0
      P[ 998] <= 9'b110000000; // Load the target box with 0
      P[ 999] <= 9'b111001001; // label: Create and set a label
      P[1000] <= 9'b001111111; // Load the constant box with 127
      P[1001] <= 9'b101000001; // Load the source box with 1
      P[1002] <= 9'b110000000; // Load the target box with 0
      P[1003] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[1004] <= 9'b011111101; // Load the constant box with 253
      P[1005] <= 9'b101000011; // Load the source box with 3
      P[1006] <= 9'b110000000; // Load the target box with 0
      P[1007] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1008] <= 9'b000010000; // Load the constant box with 16
      P[1009] <= 9'b101000011; // Load the source box with 3
      P[1010] <= 9'b110000000; // Load the target box with 0
      P[1011] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[1012] <= 9'b011111101; // Load the constant box with 253
      P[1013] <= 9'b101000011; // Load the source box with 3
      P[1014] <= 9'b110000000; // Load the target box with 0
      P[1015] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[1016] <= 9'b000001001; // Load the constant box with 9
      P[1017] <= 9'b101000000; // Load the source box with 0
      P[1018] <= 9'b110000000; // Load the target box with 0
      P[1019] <= 9'b111001001; // label: Set a label
      P[1020] <= 9'b000000000; // Load the constant box with 0
      P[1021] <= 9'b101000000; // Load the source box with 0
      P[1022] <= 9'b110000001; // Load the target box with 1
      P[1023] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[1024] <= 9'b000000111; // Load the constant box with 7
      P[1025] <= 9'b101000010; // Load the source box with 2
      P[1026] <= 9'b110000000; // Load the target box with 0
      P[1027] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[1028] <= 9'b000000000; // Load the constant box with 0
      P[1029] <= 9'b101000010; // Load the source box with 2
      P[1030] <= 9'b110000001; // Load the target box with 1
      P[1031] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[1032] <= 9'b000001101; // Load the constant box with 13
      P[1033] <= 9'b101000000; // Load the source box with 0
      P[1034] <= 9'b110000000; // Load the target box with 0
      P[1035] <= 9'b111001001; // label: Create and set a label
      P[1036] <= 9'b010000100; // Load the constant box with 132
      P[1037] <= 9'b101000001; // Load the source box with 1
      P[1038] <= 9'b110000000; // Load the target box with 0
      P[1039] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[1040] <= 9'b011111101; // Load the constant box with 253
      P[1041] <= 9'b101000011; // Load the source box with 3
      P[1042] <= 9'b110000000; // Load the target box with 0
      P[1043] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1044] <= 9'b000001000; // Load the constant box with 8
      P[1045] <= 9'b101000011; // Load the source box with 3
      P[1046] <= 9'b110000000; // Load the target box with 0
      P[1047] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[1048] <= 9'b011111101; // Load the constant box with 253
      P[1049] <= 9'b101000011; // Load the source box with 3
      P[1050] <= 9'b110000000; // Load the target box with 0
      P[1051] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[1052] <= 9'b000001010; // Load the constant box with 10
      P[1053] <= 9'b101000000; // Load the source box with 0
      P[1054] <= 9'b110000000; // Load the target box with 0
      P[1055] <= 9'b111001001; // label: Set a label
      P[1056] <= 9'b000000000; // Load the constant box with 0
      P[1057] <= 9'b101000000; // Load the source box with 0
      P[1058] <= 9'b110000001; // Load the target box with 1
      P[1059] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[1060] <= 9'b000010110; // Load the constant box with 22
      P[1061] <= 9'b101000010; // Load the source box with 2
      P[1062] <= 9'b110000000; // Load the target box with 0
      P[1063] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[1064] <= 9'b000000000; // Load the constant box with 0
      P[1065] <= 9'b101000010; // Load the source box with 2
      P[1066] <= 9'b110000001; // Load the target box with 1
      P[1067] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[1068] <= 9'b000001101; // Load the constant box with 13
      P[1069] <= 9'b101000000; // Load the source box with 0
      P[1070] <= 9'b110000000; // Load the target box with 0
      P[1071] <= 9'b111001001; // label: Create and set a label
      P[1072] <= 9'b010001000; // Load the constant box with 136
      P[1073] <= 9'b101000001; // Load the source box with 1
      P[1074] <= 9'b110000000; // Load the target box with 0
      P[1075] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[1076] <= 9'b011111101; // Load the constant box with 253
      P[1077] <= 9'b101000011; // Load the source box with 3
      P[1078] <= 9'b110000000; // Load the target box with 0
      P[1079] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1080] <= 9'b000000100; // Load the constant box with 4
      P[1081] <= 9'b101000011; // Load the source box with 3
      P[1082] <= 9'b110000000; // Load the target box with 0
      P[1083] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[1084] <= 9'b011111101; // Load the constant box with 253
      P[1085] <= 9'b101000011; // Load the source box with 3
      P[1086] <= 9'b110000000; // Load the target box with 0
      P[1087] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[1088] <= 9'b000001011; // Load the constant box with 11
      P[1089] <= 9'b101000000; // Load the source box with 0
      P[1090] <= 9'b110000000; // Load the target box with 0
      P[1091] <= 9'b111001001; // label: Set a label
      P[1092] <= 9'b000000000; // Load the constant box with 0
      P[1093] <= 9'b101000000; // Load the source box with 0
      P[1094] <= 9'b110000001; // Load the target box with 1
      P[1095] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[1096] <= 9'b000010101; // Load the constant box with 21
      P[1097] <= 9'b101000010; // Load the source box with 2
      P[1098] <= 9'b110000000; // Load the target box with 0
      P[1099] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[1100] <= 9'b000000000; // Load the constant box with 0
      P[1101] <= 9'b101000010; // Load the source box with 2
      P[1102] <= 9'b110000001; // Load the target box with 1
      P[1103] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[1104] <= 9'b000001101; // Load the constant box with 13
      P[1105] <= 9'b101000000; // Load the source box with 0
      P[1106] <= 9'b110000000; // Load the target box with 0
      P[1107] <= 9'b111001001; // label: Create and set a label
      P[1108] <= 9'b010001101; // Load the constant box with 141
      P[1109] <= 9'b101000001; // Load the source box with 1
      P[1110] <= 9'b110000000; // Load the target box with 0
      P[1111] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[1112] <= 9'b011111101; // Load the constant box with 253
      P[1113] <= 9'b101000011; // Load the source box with 3
      P[1114] <= 9'b110000000; // Load the target box with 0
      P[1115] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1116] <= 9'b000000010; // Load the constant box with 2
      P[1117] <= 9'b101000011; // Load the source box with 3
      P[1118] <= 9'b110000000; // Load the target box with 0
      P[1119] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[1120] <= 9'b011111101; // Load the constant box with 253
      P[1121] <= 9'b101000011; // Load the source box with 3
      P[1122] <= 9'b110000000; // Load the target box with 0
      P[1123] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[1124] <= 9'b000001100; // Load the constant box with 12
      P[1125] <= 9'b101000000; // Load the source box with 0
      P[1126] <= 9'b110000000; // Load the target box with 0
      P[1127] <= 9'b111001001; // label: Set a label
      P[1128] <= 9'b000000000; // Load the constant box with 0
      P[1129] <= 9'b101000000; // Load the source box with 0
      P[1130] <= 9'b110000001; // Load the target box with 1
      P[1131] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[1132] <= 9'b000010011; // Load the constant box with 19
      P[1133] <= 9'b101000010; // Load the source box with 2
      P[1134] <= 9'b110000000; // Load the target box with 0
      P[1135] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[1136] <= 9'b000000000; // Load the constant box with 0
      P[1137] <= 9'b101000010; // Load the source box with 2
      P[1138] <= 9'b110000001; // Load the target box with 1
      P[1139] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[1140] <= 9'b000001101; // Load the constant box with 13
      P[1141] <= 9'b101000000; // Load the source box with 0
      P[1142] <= 9'b110000000; // Load the target box with 0
      P[1143] <= 9'b111001001; // label: Create and set a label
      P[1144] <= 9'b010010001; // Load the constant box with 145
      P[1145] <= 9'b101000001; // Load the source box with 1
      P[1146] <= 9'b110000000; // Load the target box with 0
      P[1147] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[1148] <= 9'b011111101; // Load the constant box with 253
      P[1149] <= 9'b101000011; // Load the source box with 3
      P[1150] <= 9'b110000000; // Load the target box with 0
      P[1151] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1152] <= 9'b000000001; // Load the constant box with 1
      P[1153] <= 9'b101000011; // Load the source box with 3
      P[1154] <= 9'b110000000; // Load the target box with 0
      P[1155] <= 9'b111010101; // xor: Xor a constant with a register and save the result in the register
      P[1156] <= 9'b011111101; // Load the constant box with 253
      P[1157] <= 9'b101000011; // Load the source box with 3
      P[1158] <= 9'b110000000; // Load the target box with 0
      P[1159] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[1160] <= 9'b000001101; // Load the constant box with 13
      P[1161] <= 9'b101000000; // Load the source box with 0
      P[1162] <= 9'b110000000; // Load the target box with 0
      P[1163] <= 9'b111001001; // label: Set a label
      P[1164] <= 9'b000000010; // Load the constant box with 2
      P[1165] <= 9'b101000000; // Load the source box with 0
      P[1166] <= 9'b110000000; // Load the target box with 0
      P[1167] <= 9'b111001001; // label: Set a label
      P[1168] <= 9'b011111111; // Load the constant box with 255
      P[1169] <= 9'b101000000; // Load the source box with 0
      P[1170] <= 9'b110000000; // Load the target box with 0
      P[1171] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1172] <= 9'b011111110; // Load the constant box with 254
      P[1173] <= 9'b101000011; // Load the source box with 3
      P[1174] <= 9'b110000000; // Load the target box with 0
      P[1175] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1176] <= 9'b011111101; // Load the constant box with 253
      P[1177] <= 9'b101000100; // Load the source box with 4
      P[1178] <= 9'b110000000; // Load the target box with 0
      P[1179] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[1180] <= 9'b000011110; // Load the constant box with 30
      P[1181] <= 9'b101000101; // Load the source box with 5
      P[1182] <= 9'b110000000; // Load the target box with 0
      P[1183] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[1184] <= 9'b000000000; // Load the constant box with 0
      P[1185] <= 9'b101000000; // Load the source box with 0
      P[1186] <= 9'b110000101; // Load the target box with 5
      P[1187] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[1188] <= 9'b000000000; // Load the constant box with 0
      P[1189] <= 9'b101000101; // Load the source box with 5
      P[1190] <= 9'b110000100; // Load the target box with 4
      P[1191] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[1192] <= 9'b000000000; // Load the constant box with 0
      P[1193] <= 9'b101000101; // Load the source box with 5
      P[1194] <= 9'b110000000; // Load the target box with 0
      P[1195] <= 9'b111000110; // inc: Increment a register by one
      P[1196] <= 9'b000000000; // Load the constant box with 0
      P[1197] <= 9'b101000101; // Load the source box with 5
      P[1198] <= 9'b110000011; // Load the target box with 3
      P[1199] <= 9'b111010011; // stri: Store the contents of the first register in the location specified by the second register
      P[1200] <= 9'b000000000; // Load the constant box with 0
      P[1201] <= 9'b101000000; // Load the source box with 0
      P[1202] <= 9'b110000101; // Load the target box with 5
      P[1203] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[1204] <= 9'b001000000; // Load the constant box with 64
      P[1205] <= 9'b101000101; // Load the source box with 5
      P[1206] <= 9'b110000000; // Load the target box with 0
      P[1207] <= 9'b111000011; // cmpGt: Compare the first register with the specified constant and place a one in the register if it is greater than the constant else zero
      P[1208] <= 9'b000000001; // Load the constant box with 1
      P[1209] <= 9'b101000101; // Load the source box with 5
      P[1210] <= 9'b110000000; // Load the target box with 0
      P[1211] <= 9'b111000111; // jumpIfNotZero: Jump backwards to the specified location in the program if the register is not zero - useful for constructing for loops
      P[1212] <= 9'b000000000; // Load the constant box with 0
      P[1213] <= 9'b101000000; // Load the source box with 0
      P[1214] <= 9'b110000000; // Load the target box with 0
      P[1215] <= 9'b111010110; // stop: Stop program execution
    end
  endtask

  task  automatic load_Program3;                                                // Program 3
    begin
      $display("Program 3");
      P[   0] <= 9'b000011111; // Load the constant box with 31
      P[   1] <= 9'b101000110; // Load the source box with 6
      P[   2] <= 9'b110000000; // Load the target box with 0
      P[   3] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[   4] <= 9'b010100000; // Load the constant box with 160
      P[   5] <= 9'b101000011; // Load the source box with 3
      P[   6] <= 9'b110000000; // Load the target box with 0
      P[   7] <= 9'b111001011; // ldrd: Load the first register from a memory location
      P[   8] <= 9'b000000011; // Load the constant box with 3
      P[   9] <= 9'b101000011; // Load the source box with 3
      P[  10] <= 9'b110000000; // Load the target box with 0
      P[  11] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  12] <= 9'b010011111; // Load the constant box with 159
      P[  13] <= 9'b101001000; // Load the source box with 8
      P[  14] <= 9'b110000000; // Load the target box with 0
      P[  15] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  16] <= 9'b000010101; // Load the constant box with 21
      P[  17] <= 9'b101000000; // Load the source box with 0
      P[  18] <= 9'b110000000; // Load the target box with 0
      P[  19] <= 9'b111001001; // label: Create and set a label
      P[  20] <= 9'b000000000; // Load the constant box with 0
      P[  21] <= 9'b101001101; // Load the source box with 13
      P[  22] <= 9'b110000000; // Load the target box with 0
      P[  23] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  24] <= 9'b000000000; // Load the constant box with 0
      P[  25] <= 9'b101000101; // Load the source box with 5
      P[  26] <= 9'b110000000; // Load the target box with 0
      P[  27] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[  28] <= 9'b000000000; // Load the constant box with 0
      P[  29] <= 9'b101001000; // Load the source box with 8
      P[  30] <= 9'b110000111; // Load the target box with 7
      P[  31] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  32] <= 9'b000000000; // Load the constant box with 0
      P[  33] <= 9'b101000111; // Load the source box with 7
      P[  34] <= 9'b110000111; // Load the target box with 7
      P[  35] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[  36] <= 9'b000000000; // Load the constant box with 0
      P[  37] <= 9'b101000111; // Load the source box with 7
      P[  38] <= 9'b110000101; // Load the target box with 5
      P[  39] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  40] <= 9'b000000000; // Load the constant box with 0
      P[  41] <= 9'b101000110; // Load the source box with 6
      P[  42] <= 9'b110000101; // Load the target box with 5
      P[  43] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[  44] <= 9'b000000000; // Load the constant box with 0
      P[  45] <= 9'b101000101; // Load the source box with 5
      P[  46] <= 9'b110001010; // Load the target box with 10
      P[  47] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  48] <= 9'b000000000; // Load the constant box with 0
      P[  49] <= 9'b101000011; // Load the source box with 3
      P[  50] <= 9'b110001010; // Load the target box with 10
      P[  51] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[  52] <= 9'b000001000; // Load the constant box with 8
      P[  53] <= 9'b101001010; // Load the source box with 10
      P[  54] <= 9'b110000000; // Load the target box with 0
      P[  55] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[  56] <= 9'b000000000; // Load the constant box with 0
      P[  57] <= 9'b101001101; // Load the source box with 13
      P[  58] <= 9'b110000000; // Load the target box with 0
      P[  59] <= 9'b111000110; // inc: Increment a register by one
      P[  60] <= 9'b000000010; // Load the constant box with 2
      P[  61] <= 9'b101000000; // Load the source box with 0
      P[  62] <= 9'b110000000; // Load the target box with 0
      P[  63] <= 9'b111001001; // label: Set a label
      P[  64] <= 9'b000000001; // Load the constant box with 1
      P[  65] <= 9'b101000111; // Load the source box with 7
      P[  66] <= 9'b110000000; // Load the target box with 0
      P[  67] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[  68] <= 9'b000000000; // Load the constant box with 0
      P[  69] <= 9'b101000111; // Load the source box with 7
      P[  70] <= 9'b110000101; // Load the target box with 5
      P[  71] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  72] <= 9'b000000000; // Load the constant box with 0
      P[  73] <= 9'b101000110; // Load the source box with 6
      P[  74] <= 9'b110000101; // Load the target box with 5
      P[  75] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[  76] <= 9'b000000000; // Load the constant box with 0
      P[  77] <= 9'b101000101; // Load the source box with 5
      P[  78] <= 9'b110001010; // Load the target box with 10
      P[  79] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[  80] <= 9'b000000000; // Load the constant box with 0
      P[  81] <= 9'b101000011; // Load the source box with 3
      P[  82] <= 9'b110001010; // Load the target box with 10
      P[  83] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[  84] <= 9'b000001100; // Load the constant box with 12
      P[  85] <= 9'b101001010; // Load the source box with 10
      P[  86] <= 9'b110000000; // Load the target box with 0
      P[  87] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[  88] <= 9'b000000000; // Load the constant box with 0
      P[  89] <= 9'b101001101; // Load the source box with 13
      P[  90] <= 9'b110000000; // Load the target box with 0
      P[  91] <= 9'b111000110; // inc: Increment a register by one
      P[  92] <= 9'b000000011; // Load the constant box with 3
      P[  93] <= 9'b101000000; // Load the source box with 0
      P[  94] <= 9'b110000000; // Load the target box with 0
      P[  95] <= 9'b111001001; // label: Set a label
      P[  96] <= 9'b000000001; // Load the constant box with 1
      P[  97] <= 9'b101000111; // Load the source box with 7
      P[  98] <= 9'b110000000; // Load the target box with 0
      P[  99] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 100] <= 9'b000000000; // Load the constant box with 0
      P[ 101] <= 9'b101000111; // Load the source box with 7
      P[ 102] <= 9'b110000101; // Load the target box with 5
      P[ 103] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 104] <= 9'b000000000; // Load the constant box with 0
      P[ 105] <= 9'b101000110; // Load the source box with 6
      P[ 106] <= 9'b110000101; // Load the target box with 5
      P[ 107] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 108] <= 9'b000000000; // Load the constant box with 0
      P[ 109] <= 9'b101000101; // Load the source box with 5
      P[ 110] <= 9'b110001010; // Load the target box with 10
      P[ 111] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 112] <= 9'b000000000; // Load the constant box with 0
      P[ 113] <= 9'b101000011; // Load the source box with 3
      P[ 114] <= 9'b110001010; // Load the target box with 10
      P[ 115] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 116] <= 9'b000010000; // Load the constant box with 16
      P[ 117] <= 9'b101001010; // Load the source box with 10
      P[ 118] <= 9'b110000000; // Load the target box with 0
      P[ 119] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 120] <= 9'b000000000; // Load the constant box with 0
      P[ 121] <= 9'b101001101; // Load the source box with 13
      P[ 122] <= 9'b110000000; // Load the target box with 0
      P[ 123] <= 9'b111000110; // inc: Increment a register by one
      P[ 124] <= 9'b000000100; // Load the constant box with 4
      P[ 125] <= 9'b101000000; // Load the source box with 0
      P[ 126] <= 9'b110000000; // Load the target box with 0
      P[ 127] <= 9'b111001001; // label: Set a label
      P[ 128] <= 9'b000000001; // Load the constant box with 1
      P[ 129] <= 9'b101000111; // Load the source box with 7
      P[ 130] <= 9'b110000000; // Load the target box with 0
      P[ 131] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 132] <= 9'b000000000; // Load the constant box with 0
      P[ 133] <= 9'b101000111; // Load the source box with 7
      P[ 134] <= 9'b110000101; // Load the target box with 5
      P[ 135] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 136] <= 9'b000000000; // Load the constant box with 0
      P[ 137] <= 9'b101000110; // Load the source box with 6
      P[ 138] <= 9'b110000101; // Load the target box with 5
      P[ 139] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 140] <= 9'b000000000; // Load the constant box with 0
      P[ 141] <= 9'b101000101; // Load the source box with 5
      P[ 142] <= 9'b110001010; // Load the target box with 10
      P[ 143] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 144] <= 9'b000000000; // Load the constant box with 0
      P[ 145] <= 9'b101000011; // Load the source box with 3
      P[ 146] <= 9'b110001010; // Load the target box with 10
      P[ 147] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 148] <= 9'b000010100; // Load the constant box with 20
      P[ 149] <= 9'b101001010; // Load the source box with 10
      P[ 150] <= 9'b110000000; // Load the target box with 0
      P[ 151] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 152] <= 9'b000000000; // Load the constant box with 0
      P[ 153] <= 9'b101001101; // Load the source box with 13
      P[ 154] <= 9'b110000000; // Load the target box with 0
      P[ 155] <= 9'b111000110; // inc: Increment a register by one
      P[ 156] <= 9'b000000101; // Load the constant box with 5
      P[ 157] <= 9'b101000000; // Load the source box with 0
      P[ 158] <= 9'b110000000; // Load the target box with 0
      P[ 159] <= 9'b111001001; // label: Set a label
      P[ 160] <= 9'b000000000; // Load the constant box with 0
      P[ 161] <= 9'b101001101; // Load the source box with 13
      P[ 162] <= 9'b110000000; // Load the target box with 0
      P[ 163] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 164] <= 9'b000010110; // Load the constant box with 22
      P[ 165] <= 9'b101001101; // Load the source box with 13
      P[ 166] <= 9'b110000000; // Load the target box with 0
      P[ 167] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 168] <= 9'b000000000; // Load the constant box with 0
      P[ 169] <= 9'b101000001; // Load the source box with 1
      P[ 170] <= 9'b110000000; // Load the target box with 0
      P[ 171] <= 9'b111000110; // inc: Increment a register by one
      P[ 172] <= 9'b000000110; // Load the constant box with 6
      P[ 173] <= 9'b101000000; // Load the source box with 0
      P[ 174] <= 9'b110000000; // Load the target box with 0
      P[ 175] <= 9'b111001001; // label: Set a label
      P[ 176] <= 9'b000000000; // Load the constant box with 0
      P[ 177] <= 9'b101001000; // Load the source box with 8
      P[ 178] <= 9'b110001001; // Load the target box with 9
      P[ 179] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 180] <= 9'b010011111; // Load the constant box with 159
      P[ 181] <= 9'b101001001; // Load the source box with 9
      P[ 182] <= 9'b110000000; // Load the target box with 0
      P[ 183] <= 9'b111000100; // cmpLt: Compare the first register with the specified constant and place a one in the register if it is less than the constant else zero
      P[ 184] <= 9'b001001100; // Load the constant box with 76
      P[ 185] <= 9'b101001001; // Load the source box with 9
      P[ 186] <= 9'b110000000; // Load the target box with 0
      P[ 187] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 188] <= 9'b000000000; // Load the constant box with 0
      P[ 189] <= 9'b101001100; // Load the source box with 12
      P[ 190] <= 9'b110000000; // Load the target box with 0
      P[ 191] <= 9'b111001010; // ldrc: Load the first register from a constant
      P[ 192] <= 9'b000000000; // Load the constant box with 0
      P[ 193] <= 9'b101001000; // Load the source box with 8
      P[ 194] <= 9'b110000100; // Load the target box with 4
      P[ 195] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 196] <= 9'b000000000; // Load the constant box with 0
      P[ 197] <= 9'b101000100; // Load the source box with 4
      P[ 198] <= 9'b110000000; // Load the target box with 0
      P[ 199] <= 9'b111000110; // inc: Increment a register by one
      P[ 200] <= 9'b000000000; // Load the constant box with 0
      P[ 201] <= 9'b101000100; // Load the source box with 4
      P[ 202] <= 9'b110000100; // Load the target box with 4
      P[ 203] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[ 204] <= 9'b000001000; // Load the constant box with 8
      P[ 205] <= 9'b101000100; // Load the source box with 4
      P[ 206] <= 9'b110000000; // Load the target box with 0
      P[ 207] <= 9'b111010000; // sl: Shift the first register left by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 208] <= 9'b000000000; // Load the constant box with 0
      P[ 209] <= 9'b101001000; // Load the source box with 8
      P[ 210] <= 9'b110000101; // Load the target box with 5
      P[ 211] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 212] <= 9'b000000000; // Load the constant box with 0
      P[ 213] <= 9'b101000101; // Load the source box with 5
      P[ 214] <= 9'b110000101; // Load the target box with 5
      P[ 215] <= 9'b111001100; // ldri: Load the first register from the memory location specified by the second register
      P[ 216] <= 9'b000000000; // Load the constant box with 0
      P[ 217] <= 9'b101000101; // Load the source box with 5
      P[ 218] <= 9'b110000100; // Load the target box with 4
      P[ 219] <= 9'b111001111; // or: Or the first and second registers together and replace the first register with the result
      P[ 220] <= 9'b000000000; // Load the constant box with 0
      P[ 221] <= 9'b101000100; // Load the source box with 4
      P[ 222] <= 9'b110000101; // Load the target box with 5
      P[ 223] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 224] <= 9'b000000000; // Load the constant box with 0
      P[ 225] <= 9'b101000110; // Load the source box with 6
      P[ 226] <= 9'b110000101; // Load the target box with 5
      P[ 227] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 228] <= 9'b000000000; // Load the constant box with 0
      P[ 229] <= 9'b101000101; // Load the source box with 5
      P[ 230] <= 9'b110001010; // Load the target box with 10
      P[ 231] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 232] <= 9'b000000000; // Load the constant box with 0
      P[ 233] <= 9'b101000011; // Load the source box with 3
      P[ 234] <= 9'b110001010; // Load the target box with 10
      P[ 235] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 236] <= 9'b000011111; // Load the constant box with 31
      P[ 237] <= 9'b101001010; // Load the source box with 10
      P[ 238] <= 9'b110000000; // Load the target box with 0
      P[ 239] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 240] <= 9'b000000000; // Load the constant box with 0
      P[ 241] <= 9'b101001100; // Load the source box with 12
      P[ 242] <= 9'b110000000; // Load the target box with 0
      P[ 243] <= 9'b111000110; // inc: Increment a register by one
      P[ 244] <= 9'b000001000; // Load the constant box with 8
      P[ 245] <= 9'b101000000; // Load the source box with 0
      P[ 246] <= 9'b110000000; // Load the target box with 0
      P[ 247] <= 9'b111001001; // label: Set a label
      P[ 248] <= 9'b000000001; // Load the constant box with 1
      P[ 249] <= 9'b101000100; // Load the source box with 4
      P[ 250] <= 9'b110000000; // Load the target box with 0
      P[ 251] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 252] <= 9'b000000000; // Load the constant box with 0
      P[ 253] <= 9'b101000100; // Load the source box with 4
      P[ 254] <= 9'b110000101; // Load the target box with 5
      P[ 255] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 256] <= 9'b000000000; // Load the constant box with 0
      P[ 257] <= 9'b101000110; // Load the source box with 6
      P[ 258] <= 9'b110000101; // Load the target box with 5
      P[ 259] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 260] <= 9'b000000000; // Load the constant box with 0
      P[ 261] <= 9'b101000101; // Load the source box with 5
      P[ 262] <= 9'b110001010; // Load the target box with 10
      P[ 263] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 264] <= 9'b000000000; // Load the constant box with 0
      P[ 265] <= 9'b101000011; // Load the source box with 3
      P[ 266] <= 9'b110001010; // Load the target box with 10
      P[ 267] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 268] <= 9'b000100011; // Load the constant box with 35
      P[ 269] <= 9'b101001010; // Load the source box with 10
      P[ 270] <= 9'b110000000; // Load the target box with 0
      P[ 271] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 272] <= 9'b000000000; // Load the constant box with 0
      P[ 273] <= 9'b101001100; // Load the source box with 12
      P[ 274] <= 9'b110000000; // Load the target box with 0
      P[ 275] <= 9'b111000110; // inc: Increment a register by one
      P[ 276] <= 9'b000001001; // Load the constant box with 9
      P[ 277] <= 9'b101000000; // Load the source box with 0
      P[ 278] <= 9'b110000000; // Load the target box with 0
      P[ 279] <= 9'b111001001; // label: Set a label
      P[ 280] <= 9'b000000001; // Load the constant box with 1
      P[ 281] <= 9'b101000100; // Load the source box with 4
      P[ 282] <= 9'b110000000; // Load the target box with 0
      P[ 283] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 284] <= 9'b000000000; // Load the constant box with 0
      P[ 285] <= 9'b101000100; // Load the source box with 4
      P[ 286] <= 9'b110000101; // Load the target box with 5
      P[ 287] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 288] <= 9'b000000000; // Load the constant box with 0
      P[ 289] <= 9'b101000110; // Load the source box with 6
      P[ 290] <= 9'b110000101; // Load the target box with 5
      P[ 291] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 292] <= 9'b000000000; // Load the constant box with 0
      P[ 293] <= 9'b101000101; // Load the source box with 5
      P[ 294] <= 9'b110001010; // Load the target box with 10
      P[ 295] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 296] <= 9'b000000000; // Load the constant box with 0
      P[ 297] <= 9'b101000011; // Load the source box with 3
      P[ 298] <= 9'b110001010; // Load the target box with 10
      P[ 299] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 300] <= 9'b000100111; // Load the constant box with 39
      P[ 301] <= 9'b101001010; // Load the source box with 10
      P[ 302] <= 9'b110000000; // Load the target box with 0
      P[ 303] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 304] <= 9'b000000000; // Load the constant box with 0
      P[ 305] <= 9'b101001100; // Load the source box with 12
      P[ 306] <= 9'b110000000; // Load the target box with 0
      P[ 307] <= 9'b111000110; // inc: Increment a register by one
      P[ 308] <= 9'b000001010; // Load the constant box with 10
      P[ 309] <= 9'b101000000; // Load the source box with 0
      P[ 310] <= 9'b110000000; // Load the target box with 0
      P[ 311] <= 9'b111001001; // label: Set a label
      P[ 312] <= 9'b000000001; // Load the constant box with 1
      P[ 313] <= 9'b101000100; // Load the source box with 4
      P[ 314] <= 9'b110000000; // Load the target box with 0
      P[ 315] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 316] <= 9'b000000000; // Load the constant box with 0
      P[ 317] <= 9'b101000100; // Load the source box with 4
      P[ 318] <= 9'b110000101; // Load the target box with 5
      P[ 319] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 320] <= 9'b000000000; // Load the constant box with 0
      P[ 321] <= 9'b101000110; // Load the source box with 6
      P[ 322] <= 9'b110000101; // Load the target box with 5
      P[ 323] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 324] <= 9'b000000000; // Load the constant box with 0
      P[ 325] <= 9'b101000101; // Load the source box with 5
      P[ 326] <= 9'b110001010; // Load the target box with 10
      P[ 327] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 328] <= 9'b000000000; // Load the constant box with 0
      P[ 329] <= 9'b101000011; // Load the source box with 3
      P[ 330] <= 9'b110001010; // Load the target box with 10
      P[ 331] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 332] <= 9'b000101011; // Load the constant box with 43
      P[ 333] <= 9'b101001010; // Load the source box with 10
      P[ 334] <= 9'b110000000; // Load the target box with 0
      P[ 335] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 336] <= 9'b000000000; // Load the constant box with 0
      P[ 337] <= 9'b101001100; // Load the source box with 12
      P[ 338] <= 9'b110000000; // Load the target box with 0
      P[ 339] <= 9'b111000110; // inc: Increment a register by one
      P[ 340] <= 9'b000001011; // Load the constant box with 11
      P[ 341] <= 9'b101000000; // Load the source box with 0
      P[ 342] <= 9'b110000000; // Load the target box with 0
      P[ 343] <= 9'b111001001; // label: Set a label
      P[ 344] <= 9'b000000001; // Load the constant box with 1
      P[ 345] <= 9'b101000100; // Load the source box with 4
      P[ 346] <= 9'b110000000; // Load the target box with 0
      P[ 347] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 348] <= 9'b000000000; // Load the constant box with 0
      P[ 349] <= 9'b101000100; // Load the source box with 4
      P[ 350] <= 9'b110000101; // Load the target box with 5
      P[ 351] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 352] <= 9'b000000000; // Load the constant box with 0
      P[ 353] <= 9'b101000110; // Load the source box with 6
      P[ 354] <= 9'b110000101; // Load the target box with 5
      P[ 355] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 356] <= 9'b000000000; // Load the constant box with 0
      P[ 357] <= 9'b101000101; // Load the source box with 5
      P[ 358] <= 9'b110001010; // Load the target box with 10
      P[ 359] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 360] <= 9'b000000000; // Load the constant box with 0
      P[ 361] <= 9'b101000011; // Load the source box with 3
      P[ 362] <= 9'b110001010; // Load the target box with 10
      P[ 363] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 364] <= 9'b000101111; // Load the constant box with 47
      P[ 365] <= 9'b101001010; // Load the source box with 10
      P[ 366] <= 9'b110000000; // Load the target box with 0
      P[ 367] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 368] <= 9'b000000000; // Load the constant box with 0
      P[ 369] <= 9'b101001100; // Load the source box with 12
      P[ 370] <= 9'b110000000; // Load the target box with 0
      P[ 371] <= 9'b111000110; // inc: Increment a register by one
      P[ 372] <= 9'b000001100; // Load the constant box with 12
      P[ 373] <= 9'b101000000; // Load the source box with 0
      P[ 374] <= 9'b110000000; // Load the target box with 0
      P[ 375] <= 9'b111001001; // label: Set a label
      P[ 376] <= 9'b000000001; // Load the constant box with 1
      P[ 377] <= 9'b101000100; // Load the source box with 4
      P[ 378] <= 9'b110000000; // Load the target box with 0
      P[ 379] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 380] <= 9'b000000000; // Load the constant box with 0
      P[ 381] <= 9'b101000100; // Load the source box with 4
      P[ 382] <= 9'b110000101; // Load the target box with 5
      P[ 383] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 384] <= 9'b000000000; // Load the constant box with 0
      P[ 385] <= 9'b101000110; // Load the source box with 6
      P[ 386] <= 9'b110000101; // Load the target box with 5
      P[ 387] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 388] <= 9'b000000000; // Load the constant box with 0
      P[ 389] <= 9'b101000101; // Load the source box with 5
      P[ 390] <= 9'b110001010; // Load the target box with 10
      P[ 391] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 392] <= 9'b000000000; // Load the constant box with 0
      P[ 393] <= 9'b101000011; // Load the source box with 3
      P[ 394] <= 9'b110001010; // Load the target box with 10
      P[ 395] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 396] <= 9'b000110011; // Load the constant box with 51
      P[ 397] <= 9'b101001010; // Load the source box with 10
      P[ 398] <= 9'b110000000; // Load the target box with 0
      P[ 399] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 400] <= 9'b000000000; // Load the constant box with 0
      P[ 401] <= 9'b101001100; // Load the source box with 12
      P[ 402] <= 9'b110000000; // Load the target box with 0
      P[ 403] <= 9'b111000110; // inc: Increment a register by one
      P[ 404] <= 9'b000001101; // Load the constant box with 13
      P[ 405] <= 9'b101000000; // Load the source box with 0
      P[ 406] <= 9'b110000000; // Load the target box with 0
      P[ 407] <= 9'b111001001; // label: Set a label
      P[ 408] <= 9'b000000001; // Load the constant box with 1
      P[ 409] <= 9'b101000100; // Load the source box with 4
      P[ 410] <= 9'b110000000; // Load the target box with 0
      P[ 411] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 412] <= 9'b000000000; // Load the constant box with 0
      P[ 413] <= 9'b101000100; // Load the source box with 4
      P[ 414] <= 9'b110000101; // Load the target box with 5
      P[ 415] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 416] <= 9'b000000000; // Load the constant box with 0
      P[ 417] <= 9'b101000110; // Load the source box with 6
      P[ 418] <= 9'b110000101; // Load the target box with 5
      P[ 419] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 420] <= 9'b000000000; // Load the constant box with 0
      P[ 421] <= 9'b101000101; // Load the source box with 5
      P[ 422] <= 9'b110001010; // Load the target box with 10
      P[ 423] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 424] <= 9'b000000000; // Load the constant box with 0
      P[ 425] <= 9'b101000011; // Load the source box with 3
      P[ 426] <= 9'b110001010; // Load the target box with 10
      P[ 427] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 428] <= 9'b000110111; // Load the constant box with 55
      P[ 429] <= 9'b101001010; // Load the source box with 10
      P[ 430] <= 9'b110000000; // Load the target box with 0
      P[ 431] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 432] <= 9'b000000000; // Load the constant box with 0
      P[ 433] <= 9'b101001100; // Load the source box with 12
      P[ 434] <= 9'b110000000; // Load the target box with 0
      P[ 435] <= 9'b111000110; // inc: Increment a register by one
      P[ 436] <= 9'b000001110; // Load the constant box with 14
      P[ 437] <= 9'b101000000; // Load the source box with 0
      P[ 438] <= 9'b110000000; // Load the target box with 0
      P[ 439] <= 9'b111001001; // label: Set a label
      P[ 440] <= 9'b000000001; // Load the constant box with 1
      P[ 441] <= 9'b101000100; // Load the source box with 4
      P[ 442] <= 9'b110000000; // Load the target box with 0
      P[ 443] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 444] <= 9'b000000000; // Load the constant box with 0
      P[ 445] <= 9'b101000100; // Load the source box with 4
      P[ 446] <= 9'b110000101; // Load the target box with 5
      P[ 447] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 448] <= 9'b000000000; // Load the constant box with 0
      P[ 449] <= 9'b101000110; // Load the source box with 6
      P[ 450] <= 9'b110000101; // Load the target box with 5
      P[ 451] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 452] <= 9'b000000000; // Load the constant box with 0
      P[ 453] <= 9'b101000101; // Load the source box with 5
      P[ 454] <= 9'b110001010; // Load the target box with 10
      P[ 455] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 456] <= 9'b000000000; // Load the constant box with 0
      P[ 457] <= 9'b101000011; // Load the source box with 3
      P[ 458] <= 9'b110001010; // Load the target box with 10
      P[ 459] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 460] <= 9'b000111011; // Load the constant box with 59
      P[ 461] <= 9'b101001010; // Load the source box with 10
      P[ 462] <= 9'b110000000; // Load the target box with 0
      P[ 463] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 464] <= 9'b000000000; // Load the constant box with 0
      P[ 465] <= 9'b101001100; // Load the source box with 12
      P[ 466] <= 9'b110000000; // Load the target box with 0
      P[ 467] <= 9'b111000110; // inc: Increment a register by one
      P[ 468] <= 9'b000001111; // Load the constant box with 15
      P[ 469] <= 9'b101000000; // Load the source box with 0
      P[ 470] <= 9'b110000000; // Load the target box with 0
      P[ 471] <= 9'b111001001; // label: Set a label
      P[ 472] <= 9'b000000001; // Load the constant box with 1
      P[ 473] <= 9'b101000100; // Load the source box with 4
      P[ 474] <= 9'b110000000; // Load the target box with 0
      P[ 475] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 476] <= 9'b000000000; // Load the constant box with 0
      P[ 477] <= 9'b101000100; // Load the source box with 4
      P[ 478] <= 9'b110000101; // Load the target box with 5
      P[ 479] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 480] <= 9'b000000000; // Load the constant box with 0
      P[ 481] <= 9'b101000110; // Load the source box with 6
      P[ 482] <= 9'b110000101; // Load the target box with 5
      P[ 483] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 484] <= 9'b000000000; // Load the constant box with 0
      P[ 485] <= 9'b101000101; // Load the source box with 5
      P[ 486] <= 9'b110001010; // Load the target box with 10
      P[ 487] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 488] <= 9'b000000000; // Load the constant box with 0
      P[ 489] <= 9'b101000011; // Load the source box with 3
      P[ 490] <= 9'b110001010; // Load the target box with 10
      P[ 491] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 492] <= 9'b000111111; // Load the constant box with 63
      P[ 493] <= 9'b101001010; // Load the source box with 10
      P[ 494] <= 9'b110000000; // Load the target box with 0
      P[ 495] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 496] <= 9'b000000000; // Load the constant box with 0
      P[ 497] <= 9'b101001100; // Load the source box with 12
      P[ 498] <= 9'b110000000; // Load the target box with 0
      P[ 499] <= 9'b111000110; // inc: Increment a register by one
      P[ 500] <= 9'b000010000; // Load the constant box with 16
      P[ 501] <= 9'b101000000; // Load the source box with 0
      P[ 502] <= 9'b110000000; // Load the target box with 0
      P[ 503] <= 9'b111001001; // label: Set a label
      P[ 504] <= 9'b000000001; // Load the constant box with 1
      P[ 505] <= 9'b101000100; // Load the source box with 4
      P[ 506] <= 9'b110000000; // Load the target box with 0
      P[ 507] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 508] <= 9'b000000000; // Load the constant box with 0
      P[ 509] <= 9'b101000100; // Load the source box with 4
      P[ 510] <= 9'b110000101; // Load the target box with 5
      P[ 511] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 512] <= 9'b000000000; // Load the constant box with 0
      P[ 513] <= 9'b101000110; // Load the source box with 6
      P[ 514] <= 9'b110000101; // Load the target box with 5
      P[ 515] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 516] <= 9'b000000000; // Load the constant box with 0
      P[ 517] <= 9'b101000101; // Load the source box with 5
      P[ 518] <= 9'b110001010; // Load the target box with 10
      P[ 519] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 520] <= 9'b000000000; // Load the constant box with 0
      P[ 521] <= 9'b101000011; // Load the source box with 3
      P[ 522] <= 9'b110001010; // Load the target box with 10
      P[ 523] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 524] <= 9'b001000011; // Load the constant box with 67
      P[ 525] <= 9'b101001010; // Load the source box with 10
      P[ 526] <= 9'b110000000; // Load the target box with 0
      P[ 527] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 528] <= 9'b000000000; // Load the constant box with 0
      P[ 529] <= 9'b101001100; // Load the source box with 12
      P[ 530] <= 9'b110000000; // Load the target box with 0
      P[ 531] <= 9'b111000110; // inc: Increment a register by one
      P[ 532] <= 9'b000010001; // Load the constant box with 17
      P[ 533] <= 9'b101000000; // Load the source box with 0
      P[ 534] <= 9'b110000000; // Load the target box with 0
      P[ 535] <= 9'b111001001; // label: Set a label
      P[ 536] <= 9'b000000001; // Load the constant box with 1
      P[ 537] <= 9'b101000100; // Load the source box with 4
      P[ 538] <= 9'b110000000; // Load the target box with 0
      P[ 539] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 540] <= 9'b000000000; // Load the constant box with 0
      P[ 541] <= 9'b101000100; // Load the source box with 4
      P[ 542] <= 9'b110000101; // Load the target box with 5
      P[ 543] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 544] <= 9'b000000000; // Load the constant box with 0
      P[ 545] <= 9'b101000110; // Load the source box with 6
      P[ 546] <= 9'b110000101; // Load the target box with 5
      P[ 547] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 548] <= 9'b000000000; // Load the constant box with 0
      P[ 549] <= 9'b101000101; // Load the source box with 5
      P[ 550] <= 9'b110001010; // Load the target box with 10
      P[ 551] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 552] <= 9'b000000000; // Load the constant box with 0
      P[ 553] <= 9'b101000011; // Load the source box with 3
      P[ 554] <= 9'b110001010; // Load the target box with 10
      P[ 555] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 556] <= 9'b001000111; // Load the constant box with 71
      P[ 557] <= 9'b101001010; // Load the source box with 10
      P[ 558] <= 9'b110000000; // Load the target box with 0
      P[ 559] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 560] <= 9'b000000000; // Load the constant box with 0
      P[ 561] <= 9'b101001100; // Load the source box with 12
      P[ 562] <= 9'b110000000; // Load the target box with 0
      P[ 563] <= 9'b111000110; // inc: Increment a register by one
      P[ 564] <= 9'b000010010; // Load the constant box with 18
      P[ 565] <= 9'b101000000; // Load the source box with 0
      P[ 566] <= 9'b110000000; // Load the target box with 0
      P[ 567] <= 9'b111001001; // label: Set a label
      P[ 568] <= 9'b000000001; // Load the constant box with 1
      P[ 569] <= 9'b101000100; // Load the source box with 4
      P[ 570] <= 9'b110000000; // Load the target box with 0
      P[ 571] <= 9'b111010001; // sr: Shift the first register right by the number of bits specified by the constant filling the vacated bits with zeroes.
      P[ 572] <= 9'b000000000; // Load the constant box with 0
      P[ 573] <= 9'b101000100; // Load the source box with 4
      P[ 574] <= 9'b110000101; // Load the target box with 5
      P[ 575] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 576] <= 9'b000000000; // Load the constant box with 0
      P[ 577] <= 9'b101000110; // Load the source box with 6
      P[ 578] <= 9'b110000101; // Load the target box with 5
      P[ 579] <= 9'b111000001; // and: And the first and second registers together and replace the first register with the result
      P[ 580] <= 9'b000000000; // Load the constant box with 0
      P[ 581] <= 9'b101000101; // Load the source box with 5
      P[ 582] <= 9'b110001010; // Load the target box with 10
      P[ 583] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 584] <= 9'b000000000; // Load the constant box with 0
      P[ 585] <= 9'b101000011; // Load the source box with 3
      P[ 586] <= 9'b110001010; // Load the target box with 10
      P[ 587] <= 9'b111000010; // cmpEq: Compare two registers and set the first register to one if it is equal to the second register else zero
      P[ 588] <= 9'b001001011; // Load the constant box with 75
      P[ 589] <= 9'b101001010; // Load the source box with 10
      P[ 590] <= 9'b110000000; // Load the target box with 0
      P[ 591] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 592] <= 9'b000000000; // Load the constant box with 0
      P[ 593] <= 9'b101001100; // Load the source box with 12
      P[ 594] <= 9'b110000000; // Load the target box with 0
      P[ 595] <= 9'b111000110; // inc: Increment a register by one
      P[ 596] <= 9'b000010011; // Load the constant box with 19
      P[ 597] <= 9'b101000000; // Load the source box with 0
      P[ 598] <= 9'b110000000; // Load the target box with 0
      P[ 599] <= 9'b111001001; // label: Set a label
      P[ 600] <= 9'b000000000; // Load the constant box with 0
      P[ 601] <= 9'b101001100; // Load the source box with 12
      P[ 602] <= 9'b110000010; // Load the target box with 2
      P[ 603] <= 9'b111000000; // add: Add the first and second registers together and replace the first register with the result
      P[ 604] <= 9'b000000111; // Load the constant box with 7
      P[ 605] <= 9'b101000000; // Load the source box with 0
      P[ 606] <= 9'b110000000; // Load the target box with 0
      P[ 607] <= 9'b111001001; // label: Set a label
      P[ 608] <= 9'b000000000; // Load the constant box with 0
      P[ 609] <= 9'b101001000; // Load the source box with 8
      P[ 610] <= 9'b110001010; // Load the target box with 10
      P[ 611] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 612] <= 9'b010011111; // Load the constant box with 159
      P[ 613] <= 9'b101001010; // Load the source box with 10
      P[ 614] <= 9'b110000000; // Load the target box with 0
      P[ 615] <= 9'b111000100; // cmpLt: Compare the first register with the specified constant and place a one in the register if it is less than the constant else zero
      P[ 616] <= 9'b001010000; // Load the constant box with 80
      P[ 617] <= 9'b101001010; // Load the source box with 10
      P[ 618] <= 9'b110000000; // Load the target box with 0
      P[ 619] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 620] <= 9'b000000000; // Load the constant box with 0
      P[ 621] <= 9'b101001000; // Load the source box with 8
      P[ 622] <= 9'b110001010; // Load the target box with 10
      P[ 623] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 624] <= 9'b010000000; // Load the constant box with 128
      P[ 625] <= 9'b101001010; // Load the source box with 10
      P[ 626] <= 9'b110000000; // Load the target box with 0
      P[ 627] <= 9'b111000011; // cmpGt: Compare the first register with the specified constant and place a one in the register if it is greater than the constant else zero
      P[ 628] <= 9'b001010000; // Load the constant box with 80
      P[ 629] <= 9'b101001010; // Load the source box with 10
      P[ 630] <= 9'b110000000; // Load the target box with 0
      P[ 631] <= 9'b111001000; // jumpIfZero: Jump forwards to the specified location in the program if the register is zero - useful for constructing if statements
      P[ 632] <= 9'b000000000; // Load the constant box with 0
      P[ 633] <= 9'b101001101; // Load the source box with 13
      P[ 634] <= 9'b110000010; // Load the target box with 2
      P[ 635] <= 9'b111010100; // sub: Subtract the second register from the first register replace the first register with the result
      P[ 636] <= 9'b000010101; // Load the constant box with 21
      P[ 637] <= 9'b101000000; // Load the source box with 0
      P[ 638] <= 9'b110000000; // Load the target box with 0
      P[ 639] <= 9'b111001001; // label: Set a label
      P[ 640] <= 9'b000010100; // Load the constant box with 20
      P[ 641] <= 9'b101000000; // Load the source box with 0
      P[ 642] <= 9'b110000000; // Load the target box with 0
      P[ 643] <= 9'b111001001; // label: Set a label
      P[ 644] <= 9'b000000000; // Load the constant box with 0
      P[ 645] <= 9'b101001000; // Load the source box with 8
      P[ 646] <= 9'b110000000; // Load the target box with 0
      P[ 647] <= 9'b111000101; // dec: Decrement a register by one
      P[ 648] <= 9'b000000000; // Load the constant box with 0
      P[ 649] <= 9'b101001000; // Load the source box with 8
      P[ 650] <= 9'b110001010; // Load the target box with 10
      P[ 651] <= 9'b111001101; // ldrr: Load the first register from the second register
      P[ 652] <= 9'b001111111; // Load the constant box with 127
      P[ 653] <= 9'b101001010; // Load the source box with 10
      P[ 654] <= 9'b110000000; // Load the target box with 0
      P[ 655] <= 9'b111000011; // cmpGt: Compare the first register with the specified constant and place a one in the register if it is greater than the constant else zero
      P[ 656] <= 9'b000000010; // Load the constant box with 2
      P[ 657] <= 9'b101001010; // Load the source box with 10
      P[ 658] <= 9'b110000000; // Load the target box with 0
      P[ 659] <= 9'b111000111; // jumpIfNotZero: Jump backwards to the specified location in the program if the register is not zero - useful for constructing for loops
      P[ 660] <= 9'b011000000; // Load the constant box with 192
      P[ 661] <= 9'b101000000; // Load the source box with 0
      P[ 662] <= 9'b110000000; // Load the target box with 0
      P[ 663] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 664] <= 9'b011000001; // Load the constant box with 193
      P[ 665] <= 9'b101000001; // Load the source box with 1
      P[ 666] <= 9'b110000000; // Load the target box with 0
      P[ 667] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 668] <= 9'b011000010; // Load the constant box with 194
      P[ 669] <= 9'b101000010; // Load the source box with 2
      P[ 670] <= 9'b110000000; // Load the target box with 0
      P[ 671] <= 9'b111010010; // strd: Store the contents of the first register in the location specified by the constant
      P[ 672] <= 9'b000000000; // Load the constant box with 0
      P[ 673] <= 9'b101000000; // Load the source box with 0
      P[ 674] <= 9'b110000000; // Load the target box with 0
      P[ 675] <= 9'b111010110; // stop: Stop program execution
    end
  endtask
endmodule
