  parameter integer NInstructions = 12;

  task startTest();                                                             // MoveLong_test: load code
    begin

      code[   0] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   1] = 'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // array
      code[   2] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000001101000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   3] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000000000000000000000110100000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   4] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000001000000101010000000000000000000000000000000000000000000000000001000010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   5] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000011000000101010000000000000000000000000000000000000000000000000000011010000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   6] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000100000101010000000000000000000000000000000000000000000000000001110110000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   7] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100000000000000000000000101010000000000000000000000000000000000000000000000000000100001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   8] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100000000000000010000000101010000000000000000000000000000000000000000000000000001011001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   9] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100000000000000001000000101010000000000000000000000000000000000000000000000000000001101000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  10] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000100000000000000011000000101010000000000000000000000000000000000000000000000000001100011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[  11] = 'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000000000000000000000000000000000010000000000000001000000010101000000000000000000000000000000000000000000000000000010000000000010000000000;                                          // moveLong
    end
  endtask

  task endTest();                                                               // MoveLong_test: Evaluate results in out channel
    begin
      success = 1;
    end
  endtask
