  parameter integer NInstructions = 12;

  task startTest();                                                             // Jeq_test: load code
    begin

      code[   0] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[   1] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   2] = 'b0000000000000000000000001100010000000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // mov
      code[   3] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000101000000000000001000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000100000001000010000000000;                                          // jEq
      code[   4] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111011000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   5] = 'b0000000000000000000000001110100000000000000000000000000000000000000000000000000000000000110000000000000001000000100001000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000001000010000000000;                                          // jEq
      code[   6] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111101100000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[   7] = 'b0000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001000000000000000100000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;                                          // jmp
      code[   8] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[   9] = 'b0000000000000000000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000001011001000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // out
      code[  10] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
      code[  11] = 'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000;                                          // label
    end
  endtask

  task endTest();                                                               // Jeq_test: Evaluate results in out channel
    begin
      success = 1;
      success = success && outMem[0] == 111;
      success = success && outMem[1] == 333;
    end
  endtask
