  task startTest();                                                             // Free: load code
    begin
      NInstructionEnd = 9;

      code[   0] = 'h0000000100000000000000000000210000000000000320000000000000000000;                                                                          // array
      code[   1] = 'h0000002700000000000000000000010000000000000021000000000000000000;                                                                          // out
      code[   2] = 'h0000001400000000000000000000210000000000000320000000000000000000;                                                                          // free
      code[   3] = 'h0000000100000000000000000001210000000000000420000000000000000000;                                                                          // array
      code[   4] = 'h0000002700000000000000000000010000000000000121000000000000000000;                                                                          // out
      code[   5] = 'h0000001400000000000000000001210000000000000420000000000000000000;                                                                          // free
      code[   6] = 'h0000000100000000000000000002210000000000000520000000000000000000;                                                                          // array
      code[   7] = 'h0000002700000000000000000000010000000000000221000000000000000000;                                                                          // out
      code[   8] = 'h0000001400000000000000000002210000000000000520000000000000000000;                                                                          // free
    end
  endtask

  task endTest();                                                               // Free: Evaluate results in out channel
    begin
      success = 1;

    end
  endtask
